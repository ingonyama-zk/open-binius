module binary_tower_32b_mul (
        input ap_clk,
        input ap_rst,
        input ap_ce,
        input [31:0] a,
        input [31:0] b,
        output [31:0] ap_return
);

wire   [0:0] b0_4_fu_316_p1;
wire   [0:0] a0_212_fu_304_p1;
wire   [0:0] a1_209_fu_308_p3;
wire   [0:0] b1_120_fu_320_p3;
wire   [0:0] a_6_fu_334_p2;
wire   [0:0] b_6_fu_340_p2;
wire   [0:0] z1_fu_346_p2;
wire   [0:0] z0_fu_328_p2;
wire   [0:0] z2_fu_352_p2;
wire   [0:0] xor_ln45_fu_358_p2;
wire   [0:0] xor_ln45_1_fu_364_p2;
wire   [1:0] a1_208_fu_280_p4;
wire   [1:0] a0_211_fu_276_p1;
wire   [1:0] b1_119_fu_294_p4;
wire   [1:0] b0_3_fu_290_p1;
wire   [0:0] a0_214_fu_378_p3;
wire   [1:0] a_8_fu_386_p2;
wire   [0:0] b0_6_fu_392_p3;
wire   [1:0] b_8_fu_400_p2;
wire   [0:0] b0_5_fu_420_p2;
wire   [0:0] a0_213_fu_406_p2;
wire   [0:0] a1_210_fu_412_p3;
wire   [0:0] b1_121_fu_426_p3;
wire   [0:0] a_10_fu_440_p2;
wire   [0:0] b_10_fu_446_p2;
wire   [0:0] z1_1_fu_452_p2;
wire   [0:0] z0_2_fu_434_p2;
wire   [0:0] z2_1_fu_458_p2;
wire   [0:0] xor_ln45_2_fu_464_p2;
wire   [0:0] xor_ln45_3_fu_470_p2;
wire   [0:0] a1_211_fu_484_p3;
wire   [0:0] b1_122_fu_492_p3;
wire   [0:0] a_14_fu_506_p2;
wire   [0:0] b_14_fu_512_p2;
wire   [0:0] z1_3_fu_518_p2;
wire   [0:0] z0_3_fu_500_p2;
wire   [0:0] z2_2_fu_524_p2;
wire   [0:0] a1_9_fu_530_p2;
wire   [0:0] a0_fu_536_p2;
wire   [0:0] xor_ln28_fu_550_p2;
wire   [1:0] z1_2_fu_476_p3;
wire   [1:0] z0_1_fu_370_p3;
wire   [1:0] z2_121_fu_542_p3;
wire   [1:0] tmp_fu_556_p3;
wire   [1:0] xor_ln45_7_fu_570_p2;
wire   [1:0] xor_ln45_6_fu_564_p2;
wire   [1:0] xor_ln45_8_fu_576_p2;
wire   [1:0] xor_ln45_9_fu_582_p2;
wire   [3:0] a1_207_fu_252_p4;
wire   [3:0] a0_210_fu_248_p1;
wire   [3:0] b1_118_fu_266_p4;
wire   [3:0] b0_2_fu_262_p1;
wire   [1:0] a0_219_fu_604_p4;
wire   [3:0] a_17_fu_614_p2;
wire   [1:0] b0_11_fu_628_p4;
wire   [3:0] b_16_fu_638_p2;
wire   [0:0] a0_220_fu_596_p3;
wire   [1:0] a0_215_fu_644_p2;
wire   [0:0] b0_12_fu_620_p3;
wire   [1:0] b0_7_fu_660_p2;
wire   [0:0] b0_8_fu_690_p2;
wire   [0:0] a0_216_fu_676_p2;
wire   [0:0] a1_213_fu_682_p3;
wire   [0:0] b1_124_fu_696_p3;
wire   [0:0] a_20_fu_710_p2;
wire   [0:0] b_19_fu_716_p2;
wire   [0:0] z1_4_fu_722_p2;
wire   [0:0] z0_5_fu_704_p2;
wire   [0:0] z2_4_fu_728_p2;
wire   [0:0] xor_ln45_10_fu_734_p2;
wire   [0:0] xor_ln45_11_fu_740_p2;
wire   [1:0] a1_212_fu_650_p4;
wire   [1:0] b1_123_fu_666_p4;
wire   [0:0] a0_218_fu_754_p3;
wire   [1:0] a_22_fu_762_p2;
wire   [0:0] b0_10_fu_768_p3;
wire   [1:0] b_21_fu_776_p2;
wire   [0:0] b0_9_fu_796_p2;
wire   [0:0] a0_217_fu_782_p2;
wire   [0:0] a1_214_fu_788_p3;
wire   [0:0] b1_125_fu_802_p3;
wire   [0:0] a_24_fu_816_p2;
wire   [0:0] b_23_fu_822_p2;
wire   [0:0] z1_5_fu_828_p2;
wire   [0:0] z0_7_fu_810_p2;
wire   [0:0] z2_5_fu_834_p2;
wire   [0:0] xor_ln45_12_fu_840_p2;
wire   [0:0] xor_ln45_13_fu_846_p2;
wire   [0:0] a1_215_fu_860_p3;
wire   [0:0] b1_126_fu_868_p3;
wire   [0:0] a_28_fu_882_p2;
wire   [0:0] b_27_fu_888_p2;
wire   [0:0] z1_7_fu_894_p2;
wire   [0:0] z0_8_fu_876_p2;
wire   [0:0] z2_6_fu_900_p2;
wire   [0:0] a1_15_fu_906_p2;
wire   [0:0] a0_13_fu_912_p2;
wire   [0:0] xor_ln28_1_fu_926_p2;
wire   [1:0] z1_6_fu_852_p3;
wire   [1:0] z0_6_fu_746_p3;
wire   [1:0] z2_122_fu_918_p3;
wire   [1:0] tmp_5_fu_932_p3;
wire   [1:0] xor_ln45_17_fu_946_p2;
wire   [1:0] xor_ln45_16_fu_940_p2;
wire   [1:0] xor_ln45_18_fu_952_p2;
wire   [1:0] xor_ln45_19_fu_958_p2;
wire   [0:0] a1_217_fu_992_p3;
wire   [0:0] b1_128_fu_1000_p3;
wire   [0:0] a_34_fu_1014_p2;
wire   [0:0] b_32_fu_1020_p2;
wire   [0:0] z1_9_fu_1026_p2;
wire   [0:0] z0_9_fu_1008_p2;
wire   [0:0] z2_8_fu_1032_p2;
wire   [0:0] xor_ln45_20_fu_1038_p2;
wire   [0:0] xor_ln45_21_fu_1044_p2;
wire   [1:0] a1_216_fu_972_p4;
wire   [1:0] b1_127_fu_982_p4;
wire   [0:0] a0_222_fu_1058_p3;
wire   [1:0] a_36_fu_1066_p2;
wire   [0:0] b0_14_fu_1072_p3;
wire   [1:0] b_34_fu_1080_p2;
wire   [0:0] b0_13_fu_1100_p2;
wire   [0:0] a0_221_fu_1086_p2;
wire   [0:0] a1_218_fu_1092_p3;
wire   [0:0] b1_129_fu_1106_p3;
wire   [0:0] a_38_fu_1120_p2;
wire   [0:0] b_36_fu_1126_p2;
wire   [0:0] z1_10_fu_1132_p2;
wire   [0:0] z0_11_fu_1114_p2;
wire   [0:0] z2_9_fu_1138_p2;
wire   [0:0] xor_ln45_22_fu_1144_p2;
wire   [0:0] xor_ln45_23_fu_1150_p2;
wire   [0:0] a1_219_fu_1164_p3;
wire   [0:0] b1_130_fu_1172_p3;
wire   [0:0] a_42_fu_1186_p2;
wire   [0:0] b_40_fu_1192_p2;
wire   [0:0] z1_12_fu_1198_p2;
wire   [0:0] z0_12_fu_1180_p2;
wire   [0:0] z2_10_fu_1204_p2;
wire   [0:0] a1_21_fu_1210_p2;
wire   [0:0] a0_20_fu_1216_p2;
wire   [0:0] xor_ln28_2_fu_1230_p2;
wire   [1:0] z1_11_fu_1156_p3;
wire   [1:0] z0_10_fu_1050_p3;
wire   [1:0] z2_123_fu_1222_p3;
wire   [1:0] tmp_s_fu_1236_p3;
wire   [1:0] xor_ln45_27_fu_1250_p2;
wire   [1:0] xor_ln45_26_fu_1244_p2;
wire   [1:0] a1_220_fu_1256_p2;
wire   [1:0] a0_21_fu_1262_p2;
wire   [0:0] a0_23_fu_1276_p1;
wire   [0:0] a1_23_fu_1280_p3;
wire   [0:0] xor_ln28_3_fu_1288_p2;
wire   [1:0] tmp_1_fu_1294_p3;
wire   [1:0] xor_ln28_4_fu_1302_p2;
wire   [3:0] z1_8_fu_964_p3;
wire   [3:0] z0_4_fu_588_p3;
wire   [3:0] z2_124_fu_1268_p3;
wire   [3:0] tmp_2_fu_1308_p3;
wire   [3:0] xor_ln45_31_fu_1322_p2;
wire   [3:0] xor_ln45_30_fu_1316_p2;
wire   [3:0] xor_ln45_32_fu_1328_p2;
wire   [3:0] xor_ln45_33_fu_1334_p2;
wire   [7:0] a1_206_fu_220_p4;
wire   [7:0] a0_209_fu_212_p1;
wire   [5:0] trunc_ln43_s_fu_1376_p4;
wire   [5:0] trunc_ln38_4_fu_216_p1;
wire   [7:0] b1_117_fu_238_p4;
wire   [7:0] b0_1_fu_230_p1;
wire   [5:0] trunc_ln43_1_fu_1426_p4;
wire   [5:0] trunc_ln40_4_fu_234_p1;
wire   [3:0] a0_236_fu_1366_p4;
wire   [7:0] a_47_fu_1386_p2;
wire   [3:0] b0_28_fu_1416_p4;
wire   [7:0] b_42_fu_1436_p2;
wire   [1:0] a0_237_fu_1356_p4;
wire   [3:0] a0_223_fu_1448_p2;
wire   [1:0] b0_29_fu_1406_p4;
wire   [3:0] b0_15_fu_1464_p2;
wire   [0:0] a0_238_fu_1348_p3;
wire   [1:0] a0_224_fu_1480_p2;
wire   [0:0] b0_30_fu_1398_p3;
wire   [1:0] b0_16_fu_1496_p2;
wire   [0:0] b0_17_fu_1526_p2;
wire   [0:0] a0_225_fu_1512_p2;
wire   [0:0] a1_223_fu_1518_p3;
wire   [0:0] b1_133_fu_1532_p3;
wire   [0:0] a_51_fu_1546_p2;
wire   [0:0] b_46_fu_1552_p2;
wire   [0:0] z1_13_fu_1558_p2;
wire   [0:0] z0_14_fu_1540_p2;
wire   [0:0] z2_13_fu_1564_p2;
wire   [0:0] xor_ln45_34_fu_1570_p2;
wire   [0:0] xor_ln45_35_fu_1576_p2;
wire   [1:0] a1_222_fu_1486_p4;
wire   [1:0] b1_132_fu_1502_p4;
wire   [0:0] a0_227_fu_1590_p3;
wire   [1:0] a_53_fu_1598_p2;
wire   [0:0] b0_19_fu_1604_p3;
wire   [1:0] b_48_fu_1612_p2;
wire   [0:0] b0_18_fu_1632_p2;
wire   [0:0] a0_226_fu_1618_p2;
wire   [0:0] a1_224_fu_1624_p3;
wire   [0:0] b1_134_fu_1638_p3;
wire   [0:0] a_55_fu_1652_p2;
wire   [0:0] b_50_fu_1658_p2;
wire   [0:0] z1_14_fu_1664_p2;
wire   [0:0] z0_16_fu_1646_p2;
wire   [0:0] z2_14_fu_1670_p2;
wire   [0:0] xor_ln45_36_fu_1676_p2;
wire   [0:0] xor_ln45_37_fu_1682_p2;
wire   [0:0] a1_225_fu_1696_p3;
wire   [0:0] b1_135_fu_1704_p3;
wire   [0:0] a_59_fu_1718_p2;
wire   [0:0] b_54_fu_1724_p2;
wire   [0:0] z1_16_fu_1730_p2;
wire   [0:0] z0_17_fu_1712_p2;
wire   [0:0] z2_15_fu_1736_p2;
wire   [0:0] a1_31_fu_1742_p2;
wire   [0:0] a0_32_fu_1748_p2;
wire   [0:0] xor_ln28_5_fu_1762_p2;
wire   [1:0] z1_15_fu_1688_p3;
wire   [1:0] z0_15_fu_1582_p3;
wire   [1:0] z2_125_fu_1754_p3;
wire   [1:0] tmp_3_fu_1768_p3;
wire   [1:0] xor_ln45_41_fu_1782_p2;
wire   [1:0] xor_ln45_40_fu_1776_p2;
wire   [1:0] xor_ln45_42_fu_1788_p2;
wire   [1:0] xor_ln45_43_fu_1794_p2;
wire   [3:0] a1_221_fu_1454_p4;
wire   [3:0] b1_131_fu_1470_p4;
wire   [1:0] a0_232_fu_1816_p4;
wire   [3:0] a_62_fu_1826_p2;
wire   [1:0] b0_24_fu_1840_p4;
wire   [3:0] b_56_fu_1850_p2;
wire   [0:0] a0_233_fu_1808_p3;
wire   [1:0] a0_228_fu_1856_p2;
wire   [0:0] b0_25_fu_1832_p3;
wire   [1:0] b0_20_fu_1872_p2;
wire   [0:0] b0_21_fu_1902_p2;
wire   [0:0] a0_229_fu_1888_p2;
wire   [0:0] a1_227_fu_1894_p3;
wire   [0:0] b1_137_fu_1908_p3;
wire   [0:0] a_65_fu_1922_p2;
wire   [0:0] b_59_fu_1928_p2;
wire   [0:0] z1_17_fu_1934_p2;
wire   [0:0] z0_19_fu_1916_p2;
wire   [0:0] z2_17_fu_1940_p2;
wire   [0:0] xor_ln45_44_fu_1946_p2;
wire   [0:0] xor_ln45_45_fu_1952_p2;
wire   [1:0] a1_226_fu_1862_p4;
wire   [1:0] b1_136_fu_1878_p4;
wire   [0:0] a0_231_fu_1966_p3;
wire   [1:0] a_67_fu_1974_p2;
wire   [0:0] b0_23_fu_1980_p3;
wire   [1:0] b_61_fu_1988_p2;
wire   [0:0] b0_22_fu_2008_p2;
wire   [0:0] a0_230_fu_1994_p2;
wire   [0:0] a1_228_fu_2000_p3;
wire   [0:0] b1_138_fu_2014_p3;
wire   [0:0] a_69_fu_2028_p2;
wire   [0:0] b_63_fu_2034_p2;
wire   [0:0] z1_18_fu_2040_p2;
wire   [0:0] z0_21_fu_2022_p2;
wire   [0:0] z2_18_fu_2046_p2;
wire   [0:0] xor_ln45_46_fu_2052_p2;
wire   [0:0] xor_ln45_47_fu_2058_p2;
wire   [0:0] a1_229_fu_2072_p3;
wire   [0:0] b1_139_fu_2080_p3;
wire   [0:0] a_73_fu_2094_p2;
wire   [0:0] b_67_fu_2100_p2;
wire   [0:0] z1_20_fu_2106_p2;
wire   [0:0] z0_22_fu_2088_p2;
wire   [0:0] z2_19_fu_2112_p2;
wire   [0:0] a1_37_fu_2118_p2;
wire   [0:0] a0_39_fu_2124_p2;
wire   [0:0] xor_ln28_6_fu_2138_p2;
wire   [1:0] z1_19_fu_2064_p3;
wire   [1:0] z0_20_fu_1958_p3;
wire   [1:0] z2_126_fu_2130_p3;
wire   [1:0] tmp_4_fu_2144_p3;
wire   [1:0] xor_ln45_51_fu_2158_p2;
wire   [1:0] xor_ln45_50_fu_2152_p2;
wire   [1:0] xor_ln45_52_fu_2164_p2;
wire   [1:0] xor_ln45_53_fu_2170_p2;
wire   [5:0] xor_ln43_14_fu_1392_p2;
wire   [5:0] xor_ln33_fu_1442_p2;
wire   [0:0] a1_231_fu_2204_p3;
wire   [0:0] b1_141_fu_2212_p3;
wire   [0:0] a_79_fu_2226_p2;
wire   [0:0] b_72_fu_2232_p2;
wire   [0:0] z1_22_fu_2238_p2;
wire   [0:0] z0_23_fu_2220_p2;
wire   [0:0] z2_21_fu_2244_p2;
wire   [0:0] xor_ln45_54_fu_2250_p2;
wire   [0:0] xor_ln45_55_fu_2256_p2;
wire   [1:0] a1_230_fu_2184_p4;
wire   [1:0] b1_140_fu_2194_p4;
wire   [0:0] a0_235_fu_2270_p3;
wire   [1:0] a_81_fu_2278_p2;
wire   [0:0] b0_27_fu_2284_p3;
wire   [1:0] b_74_fu_2292_p2;
wire   [0:0] b0_26_fu_2312_p2;
wire   [0:0] a0_234_fu_2298_p2;
wire   [0:0] a1_232_fu_2304_p3;
wire   [0:0] b1_142_fu_2318_p3;
wire   [0:0] a_83_fu_2332_p2;
wire   [0:0] b_76_fu_2338_p2;
wire   [0:0] z1_23_fu_2344_p2;
wire   [0:0] z0_25_fu_2326_p2;
wire   [0:0] z2_22_fu_2350_p2;
wire   [0:0] xor_ln45_56_fu_2356_p2;
wire   [0:0] xor_ln45_57_fu_2362_p2;
wire   [0:0] a1_233_fu_2376_p3;
wire   [0:0] b1_143_fu_2384_p3;
wire   [0:0] a_87_fu_2398_p2;
wire   [0:0] b_80_fu_2404_p2;
wire   [0:0] z1_25_fu_2410_p2;
wire   [0:0] z0_26_fu_2392_p2;
wire   [0:0] z2_23_fu_2416_p2;
wire   [0:0] a1_42_fu_2422_p2;
wire   [0:0] a0_46_fu_2428_p2;
wire   [0:0] xor_ln28_7_fu_2442_p2;
wire   [1:0] z1_24_fu_2368_p3;
wire   [1:0] z0_24_fu_2262_p3;
wire   [1:0] z2_127_fu_2434_p3;
wire   [1:0] tmp_6_fu_2448_p3;
wire   [1:0] xor_ln45_61_fu_2462_p2;
wire   [1:0] xor_ln45_60_fu_2456_p2;
wire   [1:0] a1_234_fu_2468_p2;
wire   [1:0] a0_47_fu_2474_p2;
wire   [0:0] a0_48_fu_2488_p1;
wire   [0:0] a1_45_fu_2492_p3;
wire   [0:0] xor_ln28_8_fu_2500_p2;
wire   [1:0] tmp_7_fu_2506_p3;
wire   [1:0] xor_ln28_9_fu_2514_p2;
wire   [3:0] z1_21_fu_2176_p3;
wire   [3:0] z0_18_fu_1800_p3;
wire   [3:0] z2_128_fu_2480_p3;
wire   [3:0] tmp_8_fu_2520_p3;
wire   [3:0] xor_ln45_65_fu_2534_p2;
wire   [3:0] xor_ln45_64_fu_2528_p2;
wire   [3:0] xor_ln45_66_fu_2540_p2;
wire   [3:0] xor_ln45_67_fu_2546_p2;
wire   [0:0] a1_237_fu_2600_p3;
wire   [0:0] b1_146_fu_2608_p3;
wire   [0:0] a_96_fu_2622_p2;
wire   [0:0] b_86_fu_2628_p2;
wire   [0:0] z1_27_fu_2634_p2;
wire   [0:0] z0_27_fu_2616_p2;
wire   [0:0] z2_26_fu_2640_p2;
wire   [0:0] xor_ln45_68_fu_2646_p2;
wire   [0:0] xor_ln45_69_fu_2652_p2;
wire   [1:0] a1_236_fu_2580_p4;
wire   [1:0] b1_145_fu_2590_p4;
wire   [0:0] a0_240_fu_2666_p3;
wire   [1:0] a_98_fu_2674_p2;
wire   [0:0] b0_32_fu_2680_p3;
wire   [1:0] b_88_fu_2688_p2;
wire   [0:0] b0_31_fu_2708_p2;
wire   [0:0] a0_239_fu_2694_p2;
wire   [0:0] a1_238_fu_2700_p3;
wire   [0:0] b1_147_fu_2714_p3;
wire   [0:0] a_100_fu_2728_p2;
wire   [0:0] b_90_fu_2734_p2;
wire   [0:0] z1_28_fu_2740_p2;
wire   [0:0] z0_29_fu_2722_p2;
wire   [0:0] z2_27_fu_2746_p2;
wire   [0:0] xor_ln45_70_fu_2752_p2;
wire   [0:0] xor_ln45_71_fu_2758_p2;
wire   [0:0] a1_239_fu_2772_p3;
wire   [0:0] b1_148_fu_2780_p3;
wire   [0:0] a_104_fu_2794_p2;
wire   [0:0] b_94_fu_2800_p2;
wire   [0:0] z1_30_fu_2806_p2;
wire   [0:0] z0_30_fu_2788_p2;
wire   [0:0] z2_28_fu_2812_p2;
wire   [0:0] a1_52_fu_2818_p2;
wire   [0:0] a0_54_fu_2824_p2;
wire   [0:0] xor_ln28_10_fu_2838_p2;
wire   [1:0] z1_29_fu_2764_p3;
wire   [1:0] z0_28_fu_2658_p3;
wire   [1:0] z2_129_fu_2830_p3;
wire   [1:0] tmp_9_fu_2844_p3;
wire   [1:0] xor_ln45_75_fu_2858_p2;
wire   [1:0] xor_ln45_74_fu_2852_p2;
wire   [1:0] xor_ln45_76_fu_2864_p2;
wire   [1:0] xor_ln45_77_fu_2870_p2;
wire   [3:0] a1_235_fu_2560_p4;
wire   [3:0] b1_144_fu_2570_p4;
wire   [1:0] a0_245_fu_2892_p4;
wire   [3:0] a_107_fu_2902_p2;
wire   [1:0] b0_37_fu_2916_p4;
wire   [3:0] b_96_fu_2926_p2;
wire   [0:0] a0_246_fu_2884_p3;
wire   [1:0] a0_241_fu_2932_p2;
wire   [0:0] b0_38_fu_2908_p3;
wire   [1:0] b0_33_fu_2948_p2;
wire   [0:0] b0_34_fu_2978_p2;
wire   [0:0] a0_242_fu_2964_p2;
wire   [0:0] a1_241_fu_2970_p3;
wire   [0:0] b1_150_fu_2984_p3;
wire   [0:0] a_110_fu_2998_p2;
wire   [0:0] b_99_fu_3004_p2;
wire   [0:0] z1_31_fu_3010_p2;
wire   [0:0] z0_32_fu_2992_p2;
wire   [0:0] z2_30_fu_3016_p2;
wire   [0:0] xor_ln45_78_fu_3022_p2;
wire   [0:0] xor_ln45_79_fu_3028_p2;
wire   [1:0] a1_240_fu_2938_p4;
wire   [1:0] b1_149_fu_2954_p4;
wire   [0:0] a0_244_fu_3042_p3;
wire   [1:0] a_112_fu_3050_p2;
wire   [0:0] b0_36_fu_3056_p3;
wire   [1:0] b_101_fu_3064_p2;
wire   [0:0] b0_35_fu_3084_p2;
wire   [0:0] a0_243_fu_3070_p2;
wire   [0:0] a1_242_fu_3076_p3;
wire   [0:0] b1_151_fu_3090_p3;
wire   [0:0] a_114_fu_3104_p2;
wire   [0:0] b_103_fu_3110_p2;
wire   [0:0] z1_32_fu_3116_p2;
wire   [0:0] z0_34_fu_3098_p2;
wire   [0:0] z2_31_fu_3122_p2;
wire   [0:0] xor_ln45_80_fu_3128_p2;
wire   [0:0] xor_ln45_81_fu_3134_p2;
wire   [0:0] a1_243_fu_3148_p3;
wire   [0:0] b1_152_fu_3156_p3;
wire   [0:0] a_118_fu_3170_p2;
wire   [0:0] b_107_fu_3176_p2;
wire   [0:0] z1_34_fu_3182_p2;
wire   [0:0] z0_35_fu_3164_p2;
wire   [0:0] z2_32_fu_3188_p2;
wire   [0:0] a1_58_fu_3194_p2;
wire   [0:0] a0_62_fu_3200_p2;
wire   [0:0] xor_ln28_11_fu_3214_p2;
wire   [1:0] z1_33_fu_3140_p3;
wire   [1:0] z0_33_fu_3034_p3;
wire   [1:0] z2_130_fu_3206_p3;
wire   [1:0] tmp_10_fu_3220_p3;
wire   [1:0] xor_ln45_85_fu_3234_p2;
wire   [1:0] xor_ln45_84_fu_3228_p2;
wire   [1:0] xor_ln45_86_fu_3240_p2;
wire   [1:0] xor_ln45_87_fu_3246_p2;
wire   [0:0] a1_245_fu_3280_p3;
wire   [0:0] b1_154_fu_3288_p3;
wire   [0:0] a_124_fu_3302_p2;
wire   [0:0] b_112_fu_3308_p2;
wire   [0:0] z1_36_fu_3314_p2;
wire   [0:0] z0_36_fu_3296_p2;
wire   [0:0] z2_34_fu_3320_p2;
wire   [0:0] xor_ln45_88_fu_3326_p2;
wire   [0:0] xor_ln45_89_fu_3332_p2;
wire   [1:0] a1_244_fu_3260_p4;
wire   [1:0] b1_153_fu_3270_p4;
wire   [0:0] a0_248_fu_3346_p3;
wire   [1:0] a_126_fu_3354_p2;
wire   [0:0] b0_40_fu_3360_p3;
wire   [1:0] b_114_fu_3368_p2;
wire   [0:0] b0_39_fu_3388_p2;
wire   [0:0] a0_247_fu_3374_p2;
wire   [0:0] a1_246_fu_3380_p3;
wire   [0:0] b1_155_fu_3394_p3;
wire   [0:0] a_128_fu_3408_p2;
wire   [0:0] b_116_fu_3414_p2;
wire   [0:0] z1_37_fu_3420_p2;
wire   [0:0] z0_38_fu_3402_p2;
wire   [0:0] z2_35_fu_3426_p2;
wire   [0:0] xor_ln45_90_fu_3432_p2;
wire   [0:0] xor_ln45_91_fu_3438_p2;
wire   [0:0] a1_247_fu_3452_p3;
wire   [0:0] b1_156_fu_3460_p3;
wire   [0:0] a_132_fu_3474_p2;
wire   [0:0] b_120_fu_3480_p2;
wire   [0:0] z1_39_fu_3486_p2;
wire   [0:0] z0_39_fu_3468_p2;
wire   [0:0] z2_36_fu_3492_p2;
wire   [0:0] a1_63_fu_3498_p2;
wire   [0:0] a0_69_fu_3504_p2;
wire   [0:0] xor_ln28_12_fu_3518_p2;
wire   [1:0] z1_38_fu_3444_p3;
wire   [1:0] z0_37_fu_3338_p3;
wire   [1:0] z2_131_fu_3510_p3;
wire   [1:0] tmp_11_fu_3524_p3;
wire   [1:0] xor_ln45_95_fu_3538_p2;
wire   [1:0] xor_ln45_94_fu_3532_p2;
wire   [1:0] a1_248_fu_3544_p2;
wire   [1:0] a0_72_fu_3550_p2;
wire   [0:0] a0_74_fu_3564_p1;
wire   [0:0] a1_66_fu_3568_p3;
wire   [0:0] xor_ln28_13_fu_3576_p2;
wire   [1:0] tmp_12_fu_3582_p3;
wire   [1:0] xor_ln28_14_fu_3590_p2;
wire   [3:0] z1_35_fu_3252_p3;
wire   [3:0] z0_31_fu_2876_p3;
wire   [3:0] z2_132_fu_3556_p3;
wire   [3:0] tmp_13_fu_3596_p3;
wire   [3:0] xor_ln45_99_fu_3610_p2;
wire   [3:0] xor_ln45_98_fu_3604_p2;
wire   [3:0] a1_249_fu_3616_p2;
wire   [3:0] a0_75_fu_3622_p2;
wire   [0:0] a0_78_fu_3650_p3;
wire   [0:0] a1_69_fu_3658_p3;
wire   [0:0] xor_ln28_15_fu_3666_p2;
wire   [1:0] a0_76_fu_3636_p1;
wire   [1:0] tmp_14_fu_3672_p3;
wire   [1:0] xor_ln28_16_fu_3680_p2;
wire   [1:0] a1_250_fu_3640_p4;
wire   [3:0] tmp_15_fu_3686_p3;
wire   [3:0] xor_ln28_17_fu_3694_p2;
wire   [7:0] z1_26_fu_2552_p3;
wire   [7:0] z0_13_fu_1340_p3;
wire   [7:0] z2_133_fu_3628_p3;
wire   [7:0] tmp_16_fu_3700_p3;
wire   [7:0] xor_ln45_103_fu_3714_p2;
wire   [7:0] xor_ln45_102_fu_3708_p2;
wire   [7:0] xor_ln45_104_fu_3720_p2;
wire   [7:0] xor_ln45_105_fu_3726_p2;
wire   [15:0] a1_205_fu_176_p4;
wire   [15:0] a0_208_fu_160_p1;
wire   [13:0] trunc_ln43_4_fu_3798_p4;
wire   [13:0] trunc_ln38_1_fu_164_p1;
wire   [9:0] trunc_ln43_3_fu_3788_p4;
wire   [9:0] trunc_ln38_2_fu_168_p1;
wire   [11:0] trunc_ln43_2_fu_3778_p4;
wire   [11:0] trunc_ln38_3_fu_172_p1;
wire   [15:0] b1_fu_202_p4;
wire   [15:0] b0_fu_186_p1;
wire   [13:0] trunc_ln43_7_fu_3890_p4;
wire   [13:0] trunc_ln40_1_fu_190_p1;
wire   [9:0] trunc_ln43_6_fu_3880_p4;
wire   [9:0] trunc_ln40_2_fu_194_p1;
wire   [11:0] trunc_ln43_5_fu_3870_p4;
wire   [11:0] trunc_ln40_3_fu_198_p1;
wire   [7:0] a0_289_fu_3768_p4;
wire   [5:0] trunc_ln38_5_fu_3924_p4;
wire   [15:0] a_140_fu_3808_p2;
wire   [7:0] b0_81_fu_3860_p4;
wire   [5:0] trunc_ln40_5_fu_3956_p4;
wire   [15:0] b_122_fu_3900_p2;
wire   [3:0] a0_290_fu_3758_p4;
wire   [7:0] a0_249_fu_3934_p2;
wire   [3:0] b0_82_fu_3850_p4;
wire   [7:0] b0_41_fu_3966_p2;
wire   [1:0] a0_291_fu_3748_p4;
wire   [3:0] a0_250_fu_3988_p2;
wire   [1:0] b0_83_fu_3840_p4;
wire   [3:0] b0_42_fu_4004_p2;
wire   [0:0] a0_292_fu_3740_p3;
wire   [1:0] a0_251_fu_4020_p2;
wire   [0:0] b0_84_fu_3832_p3;
wire   [1:0] b0_43_fu_4036_p2;
wire   [0:0] b0_44_fu_4066_p2;
wire   [0:0] a0_252_fu_4052_p2;
wire   [0:0] a1_254_fu_4058_p3;
wire   [0:0] b1_160_fu_4072_p3;
wire   [0:0] a_145_fu_4086_p2;
wire   [0:0] b_127_fu_4092_p2;
wire   [0:0] z1_40_fu_4098_p2;
wire   [0:0] z0_41_fu_4080_p2;
wire   [0:0] z2_40_fu_4104_p2;
wire   [0:0] xor_ln45_106_fu_4110_p2;
wire   [0:0] xor_ln45_107_fu_4116_p2;
wire   [1:0] a1_253_fu_4026_p4;
wire   [1:0] b1_159_fu_4042_p4;
wire   [0:0] a0_254_fu_4130_p3;
wire   [1:0] a_147_fu_4138_p2;
wire   [0:0] b0_46_fu_4144_p3;
wire   [1:0] b_129_fu_4152_p2;
wire   [0:0] b0_45_fu_4172_p2;
wire   [0:0] a0_253_fu_4158_p2;
wire   [0:0] a1_255_fu_4164_p3;
wire   [0:0] b1_161_fu_4178_p3;
wire   [0:0] a_149_fu_4192_p2;
wire   [0:0] b_131_fu_4198_p2;
wire   [0:0] z1_41_fu_4204_p2;
wire   [0:0] z0_43_fu_4186_p2;
wire   [0:0] z2_41_fu_4210_p2;
wire   [0:0] xor_ln45_108_fu_4216_p2;
wire   [0:0] xor_ln45_109_fu_4222_p2;
wire   [0:0] a1_256_fu_4236_p3;
wire   [0:0] b1_162_fu_4244_p3;
wire   [0:0] a_153_fu_4258_p2;
wire   [0:0] b_135_fu_4264_p2;
wire   [0:0] z1_43_fu_4270_p2;
wire   [0:0] z0_44_fu_4252_p2;
wire   [0:0] z2_42_fu_4276_p2;
wire   [0:0] a1_78_fu_4282_p2;
wire   [0:0] a0_90_fu_4288_p2;
wire   [0:0] xor_ln28_18_fu_4302_p2;
wire   [1:0] z1_42_fu_4228_p3;
wire   [1:0] z0_42_fu_4122_p3;
wire   [1:0] z2_134_fu_4294_p3;
wire   [1:0] tmp_17_fu_4308_p3;
wire   [1:0] xor_ln45_113_fu_4322_p2;
wire   [1:0] xor_ln45_112_fu_4316_p2;
wire   [1:0] xor_ln45_114_fu_4328_p2;
wire   [1:0] xor_ln45_115_fu_4334_p2;
wire   [3:0] a1_252_fu_3994_p4;
wire   [3:0] b1_158_fu_4010_p4;
wire   [1:0] a0_259_fu_4356_p4;
wire   [3:0] a_156_fu_4366_p2;
wire   [1:0] b0_51_fu_4380_p4;
wire   [3:0] b_137_fu_4390_p2;
wire   [0:0] a0_260_fu_4348_p3;
wire   [1:0] a0_255_fu_4396_p2;
wire   [0:0] b0_52_fu_4372_p3;
wire   [1:0] b0_47_fu_4412_p2;
wire   [0:0] b0_48_fu_4442_p2;
wire   [0:0] a0_256_fu_4428_p2;
wire   [0:0] a1_258_fu_4434_p3;
wire   [0:0] b1_164_fu_4448_p3;
wire   [0:0] a_159_fu_4462_p2;
wire   [0:0] b_140_fu_4468_p2;
wire   [0:0] z1_44_fu_4474_p2;
wire   [0:0] z0_46_fu_4456_p2;
wire   [0:0] z2_44_fu_4480_p2;
wire   [0:0] xor_ln45_116_fu_4486_p2;
wire   [0:0] xor_ln45_117_fu_4492_p2;
wire   [1:0] a1_257_fu_4402_p4;
wire   [1:0] b1_163_fu_4418_p4;
wire   [0:0] a0_258_fu_4506_p3;
wire   [1:0] a_161_fu_4514_p2;
wire   [0:0] b0_50_fu_4520_p3;
wire   [1:0] b_142_fu_4528_p2;
wire   [0:0] b0_49_fu_4548_p2;
wire   [0:0] a0_257_fu_4534_p2;
wire   [0:0] a1_259_fu_4540_p3;
wire   [0:0] b1_165_fu_4554_p3;
wire   [0:0] a_163_fu_4568_p2;
wire   [0:0] b_144_fu_4574_p2;
wire   [0:0] z1_45_fu_4580_p2;
wire   [0:0] z0_48_fu_4562_p2;
wire   [0:0] z2_45_fu_4586_p2;
wire   [0:0] xor_ln45_118_fu_4592_p2;
wire   [0:0] xor_ln45_119_fu_4598_p2;
wire   [0:0] a1_260_fu_4612_p3;
wire   [0:0] b1_166_fu_4620_p3;
wire   [0:0] a_167_fu_4634_p2;
wire   [0:0] b_148_fu_4640_p2;
wire   [0:0] z1_47_fu_4646_p2;
wire   [0:0] z0_49_fu_4628_p2;
wire   [0:0] z2_46_fu_4652_p2;
wire   [0:0] a1_84_fu_4658_p2;
wire   [0:0] a0_97_fu_4664_p2;
wire   [0:0] xor_ln28_19_fu_4678_p2;
wire   [1:0] z1_46_fu_4604_p3;
wire   [1:0] z0_47_fu_4498_p3;
wire   [1:0] z2_135_fu_4670_p3;
wire   [1:0] tmp_18_fu_4684_p3;
wire   [1:0] xor_ln45_123_fu_4698_p2;
wire   [1:0] xor_ln45_122_fu_4692_p2;
wire   [1:0] xor_ln45_124_fu_4704_p2;
wire   [1:0] xor_ln45_125_fu_4710_p2;
wire   [5:0] xor_ln38_1_fu_3940_p2;
wire   [5:0] xor_ln40_1_fu_3972_p2;
wire   [0:0] a1_262_fu_4744_p3;
wire   [0:0] b1_168_fu_4752_p3;
wire   [0:0] a_173_fu_4766_p2;
wire   [0:0] b_153_fu_4772_p2;
wire   [0:0] z1_49_fu_4778_p2;
wire   [0:0] z0_50_fu_4760_p2;
wire   [0:0] z2_48_fu_4784_p2;
wire   [0:0] xor_ln45_126_fu_4790_p2;
wire   [0:0] xor_ln45_127_fu_4796_p2;
wire   [1:0] a1_261_fu_4724_p4;
wire   [1:0] b1_167_fu_4734_p4;
wire   [0:0] a0_262_fu_4810_p3;
wire   [1:0] a_175_fu_4818_p2;
wire   [0:0] b0_54_fu_4824_p3;
wire   [1:0] b_155_fu_4832_p2;
wire   [0:0] b0_53_fu_4852_p2;
wire   [0:0] a0_261_fu_4838_p2;
wire   [0:0] a1_263_fu_4844_p3;
wire   [0:0] b1_169_fu_4858_p3;
wire   [0:0] a_177_fu_4872_p2;
wire   [0:0] b_157_fu_4878_p2;
wire   [0:0] z1_50_fu_4884_p2;
wire   [0:0] z0_52_fu_4866_p2;
wire   [0:0] z2_49_fu_4890_p2;
wire   [0:0] xor_ln45_128_fu_4896_p2;
wire   [0:0] xor_ln45_129_fu_4902_p2;
wire   [0:0] a1_264_fu_4916_p3;
wire   [0:0] b1_170_fu_4924_p3;
wire   [0:0] a_181_fu_4938_p2;
wire   [0:0] b_161_fu_4944_p2;
wire   [0:0] z1_52_fu_4950_p2;
wire   [0:0] z0_53_fu_4932_p2;
wire   [0:0] z2_50_fu_4956_p2;
wire   [0:0] a1_90_fu_4962_p2;
wire   [0:0] a0_102_fu_4968_p2;
wire   [0:0] xor_ln28_20_fu_4982_p2;
wire   [1:0] z1_51_fu_4908_p3;
wire   [1:0] z0_51_fu_4802_p3;
wire   [1:0] z2_136_fu_4974_p3;
wire   [1:0] tmp_19_fu_4988_p3;
wire   [1:0] xor_ln45_133_fu_5002_p2;
wire   [1:0] xor_ln45_132_fu_4996_p2;
wire   [1:0] a1_265_fu_5008_p2;
wire   [1:0] a0_103_fu_5014_p2;
wire   [0:0] a0_105_fu_5028_p1;
wire   [0:0] a1_92_fu_5032_p3;
wire   [0:0] xor_ln28_21_fu_5040_p2;
wire   [1:0] tmp_20_fu_5046_p3;
wire   [1:0] xor_ln28_22_fu_5054_p2;
wire   [3:0] z1_48_fu_4716_p3;
wire   [3:0] z0_45_fu_4340_p3;
wire   [3:0] z2_137_fu_5020_p3;
wire   [3:0] tmp_21_fu_5060_p3;
wire   [3:0] xor_ln45_137_fu_5074_p2;
wire   [3:0] xor_ln45_136_fu_5068_p2;
wire   [3:0] xor_ln45_138_fu_5080_p2;
wire   [3:0] xor_ln45_139_fu_5086_p2;
wire   [7:0] a1_251_fu_3946_p4;
wire   [5:0] trunc_ln43_8_fu_5128_p4;
wire   [7:0] b1_157_fu_3978_p4;
wire   [5:0] trunc_ln43_9_fu_5178_p4;
wire   [3:0] a0_276_fu_5118_p4;
wire   [7:0] a_186_fu_5138_p2;
wire   [3:0] b0_68_fu_5168_p4;
wire   [7:0] b_163_fu_5188_p2;
wire   [1:0] a0_277_fu_5108_p4;
wire   [3:0] a0_263_fu_5200_p2;
wire   [1:0] b0_69_fu_5158_p4;
wire   [3:0] b0_55_fu_5216_p2;
wire   [0:0] a0_278_fu_5100_p3;
wire   [1:0] a0_264_fu_5232_p2;
wire   [0:0] b0_70_fu_5150_p3;
wire   [1:0] b0_56_fu_5248_p2;
wire   [0:0] b0_57_fu_5278_p2;
wire   [0:0] a0_265_fu_5264_p2;
wire   [0:0] a1_268_fu_5270_p3;
wire   [0:0] b1_173_fu_5284_p3;
wire   [0:0] a_190_fu_5298_p2;
wire   [0:0] b_167_fu_5304_p2;
wire   [0:0] z1_53_fu_5310_p2;
wire   [0:0] z0_55_fu_5292_p2;
wire   [0:0] z2_53_fu_5316_p2;
wire   [0:0] xor_ln45_140_fu_5322_p2;
wire   [0:0] xor_ln45_141_fu_5328_p2;
wire   [1:0] a1_267_fu_5238_p4;
wire   [1:0] b1_172_fu_5254_p4;
wire   [0:0] a0_267_fu_5342_p3;
wire   [1:0] a_192_fu_5350_p2;
wire   [0:0] b0_59_fu_5356_p3;
wire   [1:0] b_169_fu_5364_p2;
wire   [0:0] b0_58_fu_5384_p2;
wire   [0:0] a0_266_fu_5370_p2;
wire   [0:0] a1_269_fu_5376_p3;
wire   [0:0] b1_174_fu_5390_p3;
wire   [0:0] a_194_fu_5404_p2;
wire   [0:0] b_171_fu_5410_p2;
wire   [0:0] z1_54_fu_5416_p2;
wire   [0:0] z0_57_fu_5398_p2;
wire   [0:0] z2_54_fu_5422_p2;
wire   [0:0] xor_ln45_142_fu_5428_p2;
wire   [0:0] xor_ln45_143_fu_5434_p2;
wire   [0:0] a1_270_fu_5448_p3;
wire   [0:0] b1_175_fu_5456_p3;
wire   [0:0] a_198_fu_5470_p2;
wire   [0:0] b_175_fu_5476_p2;
wire   [0:0] z1_56_fu_5482_p2;
wire   [0:0] z0_58_fu_5464_p2;
wire   [0:0] z2_55_fu_5488_p2;
wire   [0:0] a1_99_fu_5494_p2;
wire   [0:0] a0_114_fu_5500_p2;
wire   [0:0] xor_ln28_23_fu_5514_p2;
wire   [1:0] z1_55_fu_5440_p3;
wire   [1:0] z0_56_fu_5334_p3;
wire   [1:0] z2_138_fu_5506_p3;
wire   [1:0] tmp_22_fu_5520_p3;
wire   [1:0] xor_ln45_147_fu_5534_p2;
wire   [1:0] xor_ln45_146_fu_5528_p2;
wire   [1:0] xor_ln45_148_fu_5540_p2;
wire   [1:0] xor_ln45_149_fu_5546_p2;
wire   [3:0] a1_266_fu_5206_p4;
wire   [3:0] b1_171_fu_5222_p4;
wire   [1:0] a0_272_fu_5568_p4;
wire   [3:0] a_201_fu_5578_p2;
wire   [1:0] b0_64_fu_5592_p4;
wire   [3:0] b_177_fu_5602_p2;
wire   [0:0] a0_273_fu_5560_p3;
wire   [1:0] a0_268_fu_5608_p2;
wire   [0:0] b0_65_fu_5584_p3;
wire   [1:0] b0_60_fu_5624_p2;
wire   [0:0] b0_61_fu_5654_p2;
wire   [0:0] a0_269_fu_5640_p2;
wire   [0:0] a1_272_fu_5646_p3;
wire   [0:0] b1_177_fu_5660_p3;
wire   [0:0] a_204_fu_5674_p2;
wire   [0:0] b_180_fu_5680_p2;
wire   [0:0] z1_57_fu_5686_p2;
wire   [0:0] z0_60_fu_5668_p2;
wire   [0:0] z2_57_fu_5692_p2;
wire   [0:0] xor_ln45_150_fu_5698_p2;
wire   [0:0] xor_ln45_151_fu_5704_p2;
wire   [1:0] a1_271_fu_5614_p4;
wire   [1:0] b1_176_fu_5630_p4;
wire   [0:0] a0_271_fu_5718_p3;
wire   [1:0] a_206_fu_5726_p2;
wire   [0:0] b0_63_fu_5732_p3;
wire   [1:0] b_182_fu_5740_p2;
wire   [0:0] b0_62_fu_5760_p2;
wire   [0:0] a0_270_fu_5746_p2;
wire   [0:0] a1_273_fu_5752_p3;
wire   [0:0] b1_178_fu_5766_p3;
wire   [0:0] a_208_fu_5780_p2;
wire   [0:0] b_184_fu_5786_p2;
wire   [0:0] z1_58_fu_5792_p2;
wire   [0:0] z0_62_fu_5774_p2;
wire   [0:0] z2_58_fu_5798_p2;
wire   [0:0] xor_ln45_152_fu_5804_p2;
wire   [0:0] xor_ln45_153_fu_5810_p2;
wire   [0:0] a1_274_fu_5824_p3;
wire   [0:0] b1_179_fu_5832_p3;
wire   [0:0] a_212_fu_5846_p2;
wire   [0:0] b_188_fu_5852_p2;
wire   [0:0] z1_60_fu_5858_p2;
wire   [0:0] z0_63_fu_5840_p2;
wire   [0:0] z2_59_fu_5864_p2;
wire   [0:0] a1_105_fu_5870_p2;
wire   [0:0] a0_123_fu_5876_p2;
wire   [0:0] xor_ln28_24_fu_5890_p2;
wire   [1:0] z1_59_fu_5816_p3;
wire   [1:0] z0_61_fu_5710_p3;
wire   [1:0] z2_139_fu_5882_p3;
wire   [1:0] tmp_23_fu_5896_p3;
wire   [1:0] xor_ln45_157_fu_5910_p2;
wire   [1:0] xor_ln45_156_fu_5904_p2;
wire   [1:0] xor_ln45_158_fu_5916_p2;
wire   [1:0] xor_ln45_159_fu_5922_p2;
wire   [5:0] xor_ln43_59_fu_5144_p2;
wire   [5:0] xor_ln33_4_fu_5194_p2;
wire   [0:0] a1_276_fu_5956_p3;
wire   [0:0] b1_181_fu_5964_p3;
wire   [0:0] a_218_fu_5978_p2;
wire   [0:0] b_193_fu_5984_p2;
wire   [0:0] z1_62_fu_5990_p2;
wire   [0:0] z0_64_fu_5972_p2;
wire   [0:0] z2_61_fu_5996_p2;
wire   [0:0] xor_ln45_160_fu_6002_p2;
wire   [0:0] xor_ln45_161_fu_6008_p2;
wire   [1:0] a1_275_fu_5936_p4;
wire   [1:0] b1_180_fu_5946_p4;
wire   [0:0] a0_275_fu_6022_p3;
wire   [1:0] a_220_fu_6030_p2;
wire   [0:0] b0_67_fu_6036_p3;
wire   [1:0] b_195_fu_6044_p2;
wire   [0:0] b0_66_fu_6064_p2;
wire   [0:0] a0_274_fu_6050_p2;
wire   [0:0] a1_277_fu_6056_p3;
wire   [0:0] b1_182_fu_6070_p3;
wire   [0:0] a_222_fu_6084_p2;
wire   [0:0] b_197_fu_6090_p2;
wire   [0:0] z1_63_fu_6096_p2;
wire   [0:0] z0_66_fu_6078_p2;
wire   [0:0] z2_62_fu_6102_p2;
wire   [0:0] xor_ln45_162_fu_6108_p2;
wire   [0:0] xor_ln45_163_fu_6114_p2;
wire   [0:0] a1_278_fu_6128_p3;
wire   [0:0] b1_183_fu_6136_p3;
wire   [0:0] a_226_fu_6150_p2;
wire   [0:0] b_201_fu_6156_p2;
wire   [0:0] z1_65_fu_6162_p2;
wire   [0:0] z0_67_fu_6144_p2;
wire   [0:0] z2_63_fu_6168_p2;
wire   [0:0] a1_112_fu_6174_p2;
wire   [0:0] a0_129_fu_6180_p2;
wire   [0:0] xor_ln28_25_fu_6194_p2;
wire   [1:0] z1_64_fu_6120_p3;
wire   [1:0] z0_65_fu_6014_p3;
wire   [1:0] z2_140_fu_6186_p3;
wire   [1:0] tmp_24_fu_6200_p3;
wire   [1:0] xor_ln45_167_fu_6214_p2;
wire   [1:0] xor_ln45_166_fu_6208_p2;
wire   [1:0] a1_279_fu_6220_p2;
wire   [1:0] a0_130_fu_6226_p2;
wire   [0:0] a0_131_fu_6240_p1;
wire   [0:0] a1_114_fu_6244_p3;
wire   [0:0] xor_ln28_26_fu_6252_p2;
wire   [1:0] tmp_25_fu_6258_p3;
wire   [1:0] xor_ln28_27_fu_6266_p2;
wire   [3:0] z1_61_fu_5928_p3;
wire   [3:0] z0_59_fu_5552_p3;
wire   [3:0] z2_141_fu_6232_p3;
wire   [3:0] tmp_26_fu_6272_p3;
wire   [3:0] xor_ln45_171_fu_6286_p2;
wire   [3:0] xor_ln45_170_fu_6280_p2;
wire   [3:0] xor_ln45_172_fu_6292_p2;
wire   [3:0] xor_ln45_173_fu_6298_p2;
wire   [11:0] xor_ln43_44_fu_3826_p2;
wire   [11:0] xor_ln33_3_fu_3918_p2;
wire   [9:0] xor_ln43_43_fu_3820_p2;
wire   [9:0] xor_ln33_2_fu_3912_p2;
wire   [0:0] a1_282_fu_6352_p3;
wire   [0:0] b1_186_fu_6360_p3;
wire   [0:0] a_235_fu_6374_p2;
wire   [0:0] b_207_fu_6380_p2;
wire   [0:0] z1_67_fu_6386_p2;
wire   [0:0] z0_68_fu_6368_p2;
wire   [0:0] z2_66_fu_6392_p2;
wire   [0:0] xor_ln45_174_fu_6398_p2;
wire   [0:0] xor_ln45_175_fu_6404_p2;
wire   [1:0] a1_281_fu_6332_p4;
wire   [1:0] b1_185_fu_6342_p4;
wire   [0:0] a0_280_fu_6418_p3;
wire   [1:0] a_237_fu_6426_p2;
wire   [0:0] b0_72_fu_6432_p3;
wire   [1:0] b_209_fu_6440_p2;
wire   [0:0] b0_71_fu_6460_p2;
wire   [0:0] a0_279_fu_6446_p2;
wire   [0:0] a1_283_fu_6452_p3;
wire   [0:0] b1_187_fu_6466_p3;
wire   [0:0] a_239_fu_6480_p2;
wire   [0:0] b_211_fu_6486_p2;
wire   [0:0] z1_68_fu_6492_p2;
wire   [0:0] z0_70_fu_6474_p2;
wire   [0:0] z2_67_fu_6498_p2;
wire   [0:0] xor_ln45_176_fu_6504_p2;
wire   [0:0] xor_ln45_177_fu_6510_p2;
wire   [0:0] a1_284_fu_6524_p3;
wire   [0:0] b1_188_fu_6532_p3;
wire   [0:0] a_243_fu_6546_p2;
wire   [0:0] b_215_fu_6552_p2;
wire   [0:0] z1_70_fu_6558_p2;
wire   [0:0] z0_71_fu_6540_p2;
wire   [0:0] z2_68_fu_6564_p2;
wire   [0:0] a1_120_fu_6570_p2;
wire   [0:0] a0_135_fu_6576_p2;
wire   [0:0] xor_ln28_28_fu_6590_p2;
wire   [1:0] z1_69_fu_6516_p3;
wire   [1:0] z0_69_fu_6410_p3;
wire   [1:0] z2_142_fu_6582_p3;
wire   [1:0] tmp_27_fu_6596_p3;
wire   [1:0] xor_ln45_181_fu_6610_p2;
wire   [1:0] xor_ln45_180_fu_6604_p2;
wire   [1:0] xor_ln45_182_fu_6616_p2;
wire   [1:0] xor_ln45_183_fu_6622_p2;
wire   [3:0] a1_280_fu_6312_p4;
wire   [3:0] b1_184_fu_6322_p4;
wire   [1:0] a0_285_fu_6644_p4;
wire   [3:0] a_246_fu_6654_p2;
wire   [1:0] b0_77_fu_6668_p4;
wire   [3:0] b_217_fu_6678_p2;
wire   [0:0] a0_286_fu_6636_p3;
wire   [1:0] a0_281_fu_6684_p2;
wire   [0:0] b0_78_fu_6660_p3;
wire   [1:0] b0_73_fu_6700_p2;
wire   [0:0] b0_74_fu_6730_p2;
wire   [0:0] a0_282_fu_6716_p2;
wire   [0:0] a1_286_fu_6722_p3;
wire   [0:0] b1_190_fu_6736_p3;
wire   [0:0] a_249_fu_6750_p2;
wire   [0:0] b_220_fu_6756_p2;
wire   [0:0] z1_71_fu_6762_p2;
wire   [0:0] z0_73_fu_6744_p2;
wire   [0:0] z2_70_fu_6768_p2;
wire   [0:0] xor_ln45_184_fu_6774_p2;
wire   [0:0] xor_ln45_185_fu_6780_p2;
wire   [1:0] a1_285_fu_6690_p4;
wire   [1:0] b1_189_fu_6706_p4;
wire   [0:0] a0_284_fu_6794_p3;
wire   [1:0] a_251_fu_6802_p2;
wire   [0:0] b0_76_fu_6808_p3;
wire   [1:0] b_222_fu_6816_p2;
wire   [0:0] b0_75_fu_6836_p2;
wire   [0:0] a0_283_fu_6822_p2;
wire   [0:0] a1_287_fu_6828_p3;
wire   [0:0] b1_191_fu_6842_p3;
wire   [0:0] a_253_fu_6856_p2;
wire   [0:0] b_224_fu_6862_p2;
wire   [0:0] z1_72_fu_6868_p2;
wire   [0:0] z0_75_fu_6850_p2;
wire   [0:0] z2_71_fu_6874_p2;
wire   [0:0] xor_ln45_186_fu_6880_p2;
wire   [0:0] xor_ln45_187_fu_6886_p2;
wire   [0:0] a1_288_fu_6900_p3;
wire   [0:0] b1_192_fu_6908_p3;
wire   [0:0] a_257_fu_6922_p2;
wire   [0:0] b_228_fu_6928_p2;
wire   [0:0] z1_74_fu_6934_p2;
wire   [0:0] z0_76_fu_6916_p2;
wire   [0:0] z2_72_fu_6940_p2;
wire   [0:0] a1_126_fu_6946_p2;
wire   [0:0] a0_140_fu_6952_p2;
wire   [0:0] xor_ln28_29_fu_6966_p2;
wire   [1:0] z1_73_fu_6892_p3;
wire   [1:0] z0_74_fu_6786_p3;
wire   [1:0] z2_143_fu_6958_p3;
wire   [1:0] tmp_28_fu_6972_p3;
wire   [1:0] xor_ln45_191_fu_6986_p2;
wire   [1:0] xor_ln45_190_fu_6980_p2;
wire   [1:0] xor_ln45_192_fu_6992_p2;
wire   [1:0] xor_ln45_193_fu_6998_p2;
wire   [13:0] xor_ln43_42_fu_3814_p2;
wire   [13:0] xor_ln33_1_fu_3906_p2;
wire   [0:0] a1_290_fu_7032_p3;
wire   [0:0] b1_194_fu_7040_p3;
wire   [0:0] a_263_fu_7054_p2;
wire   [0:0] b_233_fu_7060_p2;
wire   [0:0] z1_76_fu_7066_p2;
wire   [0:0] z0_77_fu_7048_p2;
wire   [0:0] z2_74_fu_7072_p2;
wire   [0:0] xor_ln45_194_fu_7078_p2;
wire   [0:0] xor_ln45_195_fu_7084_p2;
wire   [1:0] a1_289_fu_7012_p4;
wire   [1:0] b1_193_fu_7022_p4;
wire   [0:0] a0_288_fu_7098_p3;
wire   [1:0] a_265_fu_7106_p2;
wire   [0:0] b0_80_fu_7112_p3;
wire   [1:0] b_235_fu_7120_p2;
wire   [0:0] b0_79_fu_7140_p2;
wire   [0:0] a0_287_fu_7126_p2;
wire   [0:0] a1_291_fu_7132_p3;
wire   [0:0] b1_195_fu_7146_p3;
wire   [0:0] a_267_fu_7160_p2;
wire   [0:0] b_237_fu_7166_p2;
wire   [0:0] z1_77_fu_7172_p2;
wire   [0:0] z0_79_fu_7154_p2;
wire   [0:0] z2_75_fu_7178_p2;
wire   [0:0] xor_ln45_196_fu_7184_p2;
wire   [0:0] xor_ln45_197_fu_7190_p2;
wire   [0:0] a1_292_fu_7204_p3;
wire   [0:0] b1_196_fu_7212_p3;
wire   [0:0] a_271_fu_7226_p2;
wire   [0:0] b_241_fu_7232_p2;
wire   [0:0] z1_79_fu_7238_p2;
wire   [0:0] z0_80_fu_7220_p2;
wire   [0:0] z2_76_fu_7244_p2;
wire   [0:0] a1_133_fu_7250_p2;
wire   [0:0] a0_144_fu_7256_p2;
wire   [0:0] xor_ln28_30_fu_7270_p2;
wire   [1:0] z1_78_fu_7196_p3;
wire   [1:0] z0_78_fu_7090_p3;
wire   [1:0] z2_144_fu_7262_p3;
wire   [1:0] tmp_29_fu_7276_p3;
wire   [1:0] xor_ln45_201_fu_7290_p2;
wire   [1:0] xor_ln45_200_fu_7284_p2;
wire   [1:0] a1_293_fu_7296_p2;
wire   [1:0] a0_145_fu_7302_p2;
wire   [0:0] a0_146_fu_7316_p1;
wire   [0:0] a1_135_fu_7320_p3;
wire   [0:0] xor_ln28_31_fu_7328_p2;
wire   [1:0] tmp_30_fu_7334_p3;
wire   [1:0] xor_ln28_32_fu_7342_p2;
wire   [3:0] z1_75_fu_7004_p3;
wire   [3:0] z0_72_fu_6628_p3;
wire   [3:0] z2_145_fu_7308_p3;
wire   [3:0] tmp_31_fu_7348_p3;
wire   [3:0] xor_ln45_205_fu_7362_p2;
wire   [3:0] xor_ln45_204_fu_7356_p2;
wire   [3:0] a1_294_fu_7368_p2;
wire   [3:0] a0_147_fu_7374_p2;
wire   [0:0] a0_149_fu_7402_p3;
wire   [0:0] a1_138_fu_7410_p3;
wire   [0:0] xor_ln28_33_fu_7418_p2;
wire   [1:0] a0_148_fu_7388_p1;
wire   [1:0] tmp_32_fu_7424_p3;
wire   [1:0] xor_ln28_34_fu_7432_p2;
wire   [1:0] a1_295_fu_7392_p4;
wire   [3:0] tmp_33_fu_7438_p3;
wire   [3:0] xor_ln28_35_fu_7446_p2;
wire   [7:0] z1_66_fu_6304_p3;
wire   [7:0] z0_54_fu_5092_p3;
wire   [7:0] z2_146_fu_7380_p3;
wire   [7:0] tmp_34_fu_7452_p3;
wire   [7:0] xor_ln45_209_fu_7466_p2;
wire   [7:0] xor_ln45_208_fu_7460_p2;
wire   [7:0] xor_ln45_210_fu_7472_p2;
wire   [7:0] xor_ln45_211_fu_7478_p2;
wire   [0:0] a1_299_fu_7552_p3;
wire   [0:0] b1_200_fu_7560_p3;
wire   [0:0] a_284_fu_7574_p2;
wire   [0:0] b_248_fu_7580_p2;
wire   [0:0] z1_81_fu_7586_p2;
wire   [0:0] z0_81_fu_7568_p2;
wire   [0:0] z2_80_fu_7592_p2;
wire   [0:0] xor_ln45_212_fu_7598_p2;
wire   [0:0] xor_ln45_213_fu_7604_p2;
wire   [1:0] a1_298_fu_7532_p4;
wire   [1:0] b1_199_fu_7542_p4;
wire   [0:0] a0_294_fu_7618_p3;
wire   [1:0] a_286_fu_7626_p2;
wire   [0:0] b0_86_fu_7632_p3;
wire   [1:0] b_250_fu_7640_p2;
wire   [0:0] b0_85_fu_7660_p2;
wire   [0:0] a0_293_fu_7646_p2;
wire   [0:0] a1_300_fu_7652_p3;
wire   [0:0] b1_201_fu_7666_p3;
wire   [0:0] a_288_fu_7680_p2;
wire   [0:0] b_252_fu_7686_p2;
wire   [0:0] z1_82_fu_7692_p2;
wire   [0:0] z0_83_fu_7674_p2;
wire   [0:0] z2_81_fu_7698_p2;
wire   [0:0] xor_ln45_214_fu_7704_p2;
wire   [0:0] xor_ln45_215_fu_7710_p2;
wire   [0:0] a1_301_fu_7724_p3;
wire   [0:0] b1_202_fu_7732_p3;
wire   [0:0] a_292_fu_7746_p2;
wire   [0:0] b_256_fu_7752_p2;
wire   [0:0] z1_84_fu_7758_p2;
wire   [0:0] z0_84_fu_7740_p2;
wire   [0:0] z2_82_fu_7764_p2;
wire   [0:0] a1_147_fu_7770_p2;
wire   [0:0] a0_154_fu_7776_p2;
wire   [0:0] xor_ln28_36_fu_7790_p2;
wire   [1:0] z1_83_fu_7716_p3;
wire   [1:0] z0_82_fu_7610_p3;
wire   [1:0] z2_147_fu_7782_p3;
wire   [1:0] tmp_35_fu_7796_p3;
wire   [1:0] xor_ln45_219_fu_7810_p2;
wire   [1:0] xor_ln45_218_fu_7804_p2;
wire   [1:0] xor_ln45_220_fu_7816_p2;
wire   [1:0] xor_ln45_221_fu_7822_p2;
wire   [3:0] a1_297_fu_7512_p4;
wire   [3:0] b1_198_fu_7522_p4;
wire   [1:0] a0_299_fu_7844_p4;
wire   [3:0] a_295_fu_7854_p2;
wire   [1:0] b0_91_fu_7868_p4;
wire   [3:0] b_258_fu_7878_p2;
wire   [0:0] a0_300_fu_7836_p3;
wire   [1:0] a0_295_fu_7884_p2;
wire   [0:0] b0_92_fu_7860_p3;
wire   [1:0] b0_87_fu_7900_p2;
wire   [0:0] b0_88_fu_7930_p2;
wire   [0:0] a0_296_fu_7916_p2;
wire   [0:0] a1_303_fu_7922_p3;
wire   [0:0] b1_204_fu_7936_p3;
wire   [0:0] a_298_fu_7950_p2;
wire   [0:0] b_261_fu_7956_p2;
wire   [0:0] z1_85_fu_7962_p2;
wire   [0:0] z0_86_fu_7944_p2;
wire   [0:0] z2_84_fu_7968_p2;
wire   [0:0] xor_ln45_222_fu_7974_p2;
wire   [0:0] xor_ln45_223_fu_7980_p2;
wire   [1:0] a1_302_fu_7890_p4;
wire   [1:0] b1_203_fu_7906_p4;
wire   [0:0] a0_298_fu_7994_p3;
wire   [1:0] a_300_fu_8002_p2;
wire   [0:0] b0_90_fu_8008_p3;
wire   [1:0] b_263_fu_8016_p2;
wire   [0:0] b0_89_fu_8036_p2;
wire   [0:0] a0_297_fu_8022_p2;
wire   [0:0] a1_304_fu_8028_p3;
wire   [0:0] b1_205_fu_8042_p3;
wire   [0:0] a_302_fu_8056_p2;
wire   [0:0] b_265_fu_8062_p2;
wire   [0:0] z1_86_fu_8068_p2;
wire   [0:0] z0_88_fu_8050_p2;
wire   [0:0] z2_85_fu_8074_p2;
wire   [0:0] xor_ln45_224_fu_8080_p2;
wire   [0:0] xor_ln45_225_fu_8086_p2;
wire   [0:0] a1_305_fu_8100_p3;
wire   [0:0] b1_206_fu_8108_p3;
wire   [0:0] a_306_fu_8122_p2;
wire   [0:0] b_269_fu_8128_p2;
wire   [0:0] z1_88_fu_8134_p2;
wire   [0:0] z0_89_fu_8116_p2;
wire   [0:0] z2_86_fu_8140_p2;
wire   [0:0] a1_153_fu_8146_p2;
wire   [0:0] a0_159_fu_8152_p2;
wire   [0:0] xor_ln28_37_fu_8166_p2;
wire   [1:0] z1_87_fu_8092_p3;
wire   [1:0] z0_87_fu_7986_p3;
wire   [1:0] z2_148_fu_8158_p3;
wire   [1:0] tmp_36_fu_8172_p3;
wire   [1:0] xor_ln45_229_fu_8186_p2;
wire   [1:0] xor_ln45_228_fu_8180_p2;
wire   [1:0] xor_ln45_230_fu_8192_p2;
wire   [1:0] xor_ln45_231_fu_8198_p2;
wire   [0:0] a1_307_fu_8232_p3;
wire   [0:0] b1_208_fu_8240_p3;
wire   [0:0] a_312_fu_8254_p2;
wire   [0:0] b_274_fu_8260_p2;
wire   [0:0] z1_90_fu_8266_p2;
wire   [0:0] z0_90_fu_8248_p2;
wire   [0:0] z2_88_fu_8272_p2;
wire   [0:0] xor_ln45_232_fu_8278_p2;
wire   [0:0] xor_ln45_233_fu_8284_p2;
wire   [1:0] a1_306_fu_8212_p4;
wire   [1:0] b1_207_fu_8222_p4;
wire   [0:0] a0_302_fu_8298_p3;
wire   [1:0] a_314_fu_8306_p2;
wire   [0:0] b0_94_fu_8312_p3;
wire   [1:0] b_276_fu_8320_p2;
wire   [0:0] b0_93_fu_8340_p2;
wire   [0:0] a0_301_fu_8326_p2;
wire   [0:0] a1_308_fu_8332_p3;
wire   [0:0] b1_209_fu_8346_p3;
wire   [0:0] a_316_fu_8360_p2;
wire   [0:0] b_278_fu_8366_p2;
wire   [0:0] z1_91_fu_8372_p2;
wire   [0:0] z0_92_fu_8354_p2;
wire   [0:0] z2_89_fu_8378_p2;
wire   [0:0] xor_ln45_234_fu_8384_p2;
wire   [0:0] xor_ln45_235_fu_8390_p2;
wire   [0:0] a1_309_fu_8404_p3;
wire   [0:0] b1_210_fu_8412_p3;
wire   [0:0] a_320_fu_8426_p2;
wire   [0:0] b_282_fu_8432_p2;
wire   [0:0] z1_93_fu_8438_p2;
wire   [0:0] z0_93_fu_8420_p2;
wire   [0:0] z2_90_fu_8444_p2;
wire   [0:0] a1_159_fu_8450_p2;
wire   [0:0] a0_164_fu_8456_p2;
wire   [0:0] xor_ln28_38_fu_8470_p2;
wire   [1:0] z1_92_fu_8396_p3;
wire   [1:0] z0_91_fu_8290_p3;
wire   [1:0] z2_149_fu_8462_p3;
wire   [1:0] tmp_37_fu_8476_p3;
wire   [1:0] xor_ln45_239_fu_8490_p2;
wire   [1:0] xor_ln45_238_fu_8484_p2;
wire   [1:0] a1_310_fu_8496_p2;
wire   [1:0] a0_165_fu_8502_p2;
wire   [0:0] a0_166_fu_8516_p1;
wire   [0:0] a1_161_fu_8520_p3;
wire   [0:0] xor_ln28_39_fu_8528_p2;
wire   [1:0] tmp_38_fu_8534_p3;
wire   [1:0] xor_ln28_40_fu_8542_p2;
wire   [3:0] z1_89_fu_8204_p3;
wire   [3:0] z0_85_fu_7828_p3;
wire   [3:0] z2_150_fu_8508_p3;
wire   [3:0] tmp_39_fu_8548_p3;
wire   [3:0] xor_ln45_243_fu_8562_p2;
wire   [3:0] xor_ln45_242_fu_8556_p2;
wire   [3:0] xor_ln45_244_fu_8568_p2;
wire   [3:0] xor_ln45_245_fu_8574_p2;
wire   [7:0] a1_296_fu_7492_p4;
wire   [5:0] trunc_ln43_10_fu_8616_p4;
wire   [7:0] b1_197_fu_7502_p4;
wire   [5:0] trunc_ln43_11_fu_8666_p4;
wire   [3:0] a0_316_fu_8606_p4;
wire   [7:0] a_325_fu_8626_p2;
wire   [3:0] b0_108_fu_8656_p4;
wire   [7:0] b_284_fu_8676_p2;
wire   [1:0] a0_317_fu_8596_p4;
wire   [3:0] a0_303_fu_8688_p2;
wire   [1:0] b0_109_fu_8646_p4;
wire   [3:0] b0_95_fu_8704_p2;
wire   [0:0] a0_318_fu_8588_p3;
wire   [1:0] a0_304_fu_8720_p2;
wire   [0:0] b0_110_fu_8638_p3;
wire   [1:0] b0_96_fu_8736_p2;
wire   [0:0] b0_97_fu_8766_p2;
wire   [0:0] a0_305_fu_8752_p2;
wire   [0:0] a1_313_fu_8758_p3;
wire   [0:0] b1_213_fu_8772_p3;
wire   [0:0] a_329_fu_8786_p2;
wire   [0:0] b_288_fu_8792_p2;
wire   [0:0] z1_94_fu_8798_p2;
wire   [0:0] z0_95_fu_8780_p2;
wire   [0:0] z2_93_fu_8804_p2;
wire   [0:0] xor_ln45_246_fu_8810_p2;
wire   [0:0] xor_ln45_247_fu_8816_p2;
wire   [1:0] a1_312_fu_8726_p4;
wire   [1:0] b1_212_fu_8742_p4;
wire   [0:0] a0_307_fu_8830_p3;
wire   [1:0] a_331_fu_8838_p2;
wire   [0:0] b0_99_fu_8844_p3;
wire   [1:0] b_290_fu_8852_p2;
wire   [0:0] b0_98_fu_8872_p2;
wire   [0:0] a0_306_fu_8858_p2;
wire   [0:0] a1_314_fu_8864_p3;
wire   [0:0] b1_214_fu_8878_p3;
wire   [0:0] a_333_fu_8892_p2;
wire   [0:0] b_292_fu_8898_p2;
wire   [0:0] z1_95_fu_8904_p2;
wire   [0:0] z0_97_fu_8886_p2;
wire   [0:0] z2_94_fu_8910_p2;
wire   [0:0] xor_ln45_248_fu_8916_p2;
wire   [0:0] xor_ln45_249_fu_8922_p2;
wire   [0:0] a1_315_fu_8936_p3;
wire   [0:0] b1_215_fu_8944_p3;
wire   [0:0] a_337_fu_8958_p2;
wire   [0:0] b_296_fu_8964_p2;
wire   [0:0] z1_97_fu_8970_p2;
wire   [0:0] z0_98_fu_8952_p2;
wire   [0:0] z2_95_fu_8976_p2;
wire   [0:0] a1_168_fu_8982_p2;
wire   [0:0] a0_172_fu_8988_p2;
wire   [0:0] xor_ln28_41_fu_9002_p2;
wire   [1:0] z1_96_fu_8928_p3;
wire   [1:0] z0_96_fu_8822_p3;
wire   [1:0] z2_151_fu_8994_p3;
wire   [1:0] tmp_40_fu_9008_p3;
wire   [1:0] xor_ln45_253_fu_9022_p2;
wire   [1:0] xor_ln45_252_fu_9016_p2;
wire   [1:0] xor_ln45_254_fu_9028_p2;
wire   [1:0] xor_ln45_255_fu_9034_p2;
wire   [3:0] a1_311_fu_8694_p4;
wire   [3:0] b1_211_fu_8710_p4;
wire   [1:0] a0_312_fu_9056_p4;
wire   [3:0] a_340_fu_9066_p2;
wire   [1:0] b0_104_fu_9080_p4;
wire   [3:0] b_298_fu_9090_p2;
wire   [0:0] a0_313_fu_9048_p3;
wire   [1:0] a0_308_fu_9096_p2;
wire   [0:0] b0_105_fu_9072_p3;
wire   [1:0] b0_100_fu_9112_p2;
wire   [0:0] b0_101_fu_9142_p2;
wire   [0:0] a0_309_fu_9128_p2;
wire   [0:0] a1_317_fu_9134_p3;
wire   [0:0] b1_217_fu_9148_p3;
wire   [0:0] a_343_fu_9162_p2;
wire   [0:0] b_301_fu_9168_p2;
wire   [0:0] z1_98_fu_9174_p2;
wire   [0:0] z0_100_fu_9156_p2;
wire   [0:0] z2_97_fu_9180_p2;
wire   [0:0] xor_ln45_256_fu_9186_p2;
wire   [0:0] xor_ln45_257_fu_9192_p2;
wire   [1:0] a1_316_fu_9102_p4;
wire   [1:0] b1_216_fu_9118_p4;
wire   [0:0] a0_311_fu_9206_p3;
wire   [1:0] a_345_fu_9214_p2;
wire   [0:0] b0_103_fu_9220_p3;
wire   [1:0] b_303_fu_9228_p2;
wire   [0:0] b0_102_fu_9248_p2;
wire   [0:0] a0_310_fu_9234_p2;
wire   [0:0] a1_318_fu_9240_p3;
wire   [0:0] b1_218_fu_9254_p3;
wire   [0:0] a_347_fu_9268_p2;
wire   [0:0] b_305_fu_9274_p2;
wire   [0:0] z1_99_fu_9280_p2;
wire   [0:0] z0_102_fu_9262_p2;
wire   [0:0] z2_98_fu_9286_p2;
wire   [0:0] xor_ln45_258_fu_9292_p2;
wire   [0:0] xor_ln45_259_fu_9298_p2;
wire   [0:0] a1_319_fu_9312_p3;
wire   [0:0] b1_219_fu_9320_p3;
wire   [0:0] a_351_fu_9334_p2;
wire   [0:0] b_309_fu_9340_p2;
wire   [0:0] z1_101_fu_9346_p2;
wire   [0:0] z0_103_fu_9328_p2;
wire   [0:0] z2_99_fu_9352_p2;
wire   [0:0] a1_173_fu_9358_p2;
wire   [0:0] a0_177_fu_9364_p2;
wire   [0:0] xor_ln28_42_fu_9378_p2;
wire   [1:0] z1_100_fu_9304_p3;
wire   [1:0] z0_101_fu_9198_p3;
wire   [1:0] z2_152_fu_9370_p3;
wire   [1:0] tmp_41_fu_9384_p3;
wire   [1:0] xor_ln45_263_fu_9398_p2;
wire   [1:0] xor_ln45_262_fu_9392_p2;
wire   [1:0] xor_ln45_264_fu_9404_p2;
wire   [1:0] xor_ln45_265_fu_9410_p2;
wire   [5:0] xor_ln43_100_fu_8632_p2;
wire   [5:0] xor_ln33_5_fu_8682_p2;
wire   [0:0] a1_321_fu_9444_p3;
wire   [0:0] b1_221_fu_9452_p3;
wire   [0:0] a_357_fu_9466_p2;
wire   [0:0] b_314_fu_9472_p2;
wire   [0:0] z1_103_fu_9478_p2;
wire   [0:0] z0_104_fu_9460_p2;
wire   [0:0] z2_101_fu_9484_p2;
wire   [0:0] xor_ln45_266_fu_9490_p2;
wire   [0:0] xor_ln45_267_fu_9496_p2;
wire   [1:0] a1_320_fu_9424_p4;
wire   [1:0] b1_220_fu_9434_p4;
wire   [0:0] a0_315_fu_9510_p3;
wire   [1:0] a_359_fu_9518_p2;
wire   [0:0] b0_107_fu_9524_p3;
wire   [1:0] b_316_fu_9532_p2;
wire   [0:0] b0_106_fu_9552_p2;
wire   [0:0] a0_314_fu_9538_p2;
wire   [0:0] a1_322_fu_9544_p3;
wire   [0:0] b1_222_fu_9558_p3;
wire   [0:0] a_361_fu_9572_p2;
wire   [0:0] b_318_fu_9578_p2;
wire   [0:0] z1_104_fu_9584_p2;
wire   [0:0] z0_106_fu_9566_p2;
wire   [0:0] z2_102_fu_9590_p2;
wire   [0:0] xor_ln45_268_fu_9596_p2;
wire   [0:0] xor_ln45_269_fu_9602_p2;
wire   [0:0] a1_323_fu_9616_p3;
wire   [0:0] b1_223_fu_9624_p3;
wire   [0:0] a_365_fu_9638_p2;
wire   [0:0] b_322_fu_9644_p2;
wire   [0:0] z1_106_fu_9650_p2;
wire   [0:0] z0_107_fu_9632_p2;
wire   [0:0] z2_103_fu_9656_p2;
wire   [0:0] a1_178_fu_9662_p2;
wire   [0:0] a0_181_fu_9668_p2;
wire   [0:0] xor_ln28_43_fu_9682_p2;
wire   [1:0] z1_105_fu_9608_p3;
wire   [1:0] z0_105_fu_9502_p3;
wire   [1:0] z2_153_fu_9674_p3;
wire   [1:0] tmp_42_fu_9688_p3;
wire   [1:0] xor_ln45_273_fu_9702_p2;
wire   [1:0] xor_ln45_272_fu_9696_p2;
wire   [1:0] a1_324_fu_9708_p2;
wire   [1:0] a0_182_fu_9714_p2;
wire   [0:0] a0_183_fu_9728_p1;
wire   [0:0] a1_180_fu_9732_p3;
wire   [0:0] xor_ln28_44_fu_9740_p2;
wire   [1:0] tmp_43_fu_9746_p3;
wire   [1:0] xor_ln28_45_fu_9754_p2;
wire   [3:0] z1_102_fu_9416_p3;
wire   [3:0] z0_99_fu_9040_p3;
wire   [3:0] z2_154_fu_9720_p3;
wire   [3:0] tmp_44_fu_9760_p3;
wire   [3:0] xor_ln45_277_fu_9774_p2;
wire   [3:0] xor_ln45_276_fu_9768_p2;
wire   [3:0] xor_ln45_278_fu_9780_p2;
wire   [3:0] xor_ln45_279_fu_9786_p2;
wire   [0:0] a1_327_fu_9840_p3;
wire   [0:0] b1_226_fu_9848_p3;
wire   [0:0] a_374_fu_9862_p2;
wire   [0:0] b_328_fu_9868_p2;
wire   [0:0] z1_108_fu_9874_p2;
wire   [0:0] z0_108_fu_9856_p2;
wire   [0:0] z2_106_fu_9880_p2;
wire   [0:0] xor_ln45_280_fu_9886_p2;
wire   [0:0] xor_ln45_281_fu_9892_p2;
wire   [1:0] a1_326_fu_9820_p4;
wire   [1:0] b1_225_fu_9830_p4;
wire   [0:0] a0_320_fu_9906_p3;
wire   [1:0] a_376_fu_9914_p2;
wire   [0:0] b0_112_fu_9920_p3;
wire   [1:0] b_330_fu_9928_p2;
wire   [0:0] b0_111_fu_9948_p2;
wire   [0:0] a0_319_fu_9934_p2;
wire   [0:0] a1_328_fu_9940_p3;
wire   [0:0] b1_227_fu_9954_p3;
wire   [0:0] a_378_fu_9968_p2;
wire   [0:0] b_332_fu_9974_p2;
wire   [0:0] z1_109_fu_9980_p2;
wire   [0:0] z0_110_fu_9962_p2;
wire   [0:0] z2_107_fu_9986_p2;
wire   [0:0] xor_ln45_282_fu_9992_p2;
wire   [0:0] xor_ln45_283_fu_9998_p2;
wire   [0:0] a1_329_fu_10012_p3;
wire   [0:0] b1_228_fu_10020_p3;
wire   [0:0] a_382_fu_10034_p2;
wire   [0:0] b_336_fu_10040_p2;
wire   [0:0] z1_111_fu_10046_p2;
wire   [0:0] z0_111_fu_10028_p2;
wire   [0:0] z2_108_fu_10052_p2;
wire   [0:0] a1_186_fu_10058_p2;
wire   [0:0] a0_188_fu_10064_p2;
wire   [0:0] xor_ln28_46_fu_10078_p2;
wire   [1:0] z1_110_fu_10004_p3;
wire   [1:0] z0_109_fu_9898_p3;
wire   [1:0] z2_155_fu_10070_p3;
wire   [1:0] tmp_45_fu_10084_p3;
wire   [1:0] xor_ln45_287_fu_10098_p2;
wire   [1:0] xor_ln45_286_fu_10092_p2;
wire   [1:0] xor_ln45_288_fu_10104_p2;
wire   [1:0] xor_ln45_289_fu_10110_p2;
wire   [3:0] a1_325_fu_9800_p4;
wire   [3:0] b1_224_fu_9810_p4;
wire   [1:0] a0_325_fu_10132_p4;
wire   [3:0] a_385_fu_10142_p2;
wire   [1:0] b0_117_fu_10156_p4;
wire   [3:0] b_338_fu_10166_p2;
wire   [0:0] a0_326_fu_10124_p3;
wire   [1:0] a0_321_fu_10172_p2;
wire   [0:0] b0_118_fu_10148_p3;
wire   [1:0] b0_113_fu_10188_p2;
wire   [0:0] b0_114_fu_10218_p2;
wire   [0:0] a0_322_fu_10204_p2;
wire   [0:0] a1_331_fu_10210_p3;
wire   [0:0] b1_230_fu_10224_p3;
wire   [0:0] a_388_fu_10238_p2;
wire   [0:0] b_341_fu_10244_p2;
wire   [0:0] z1_112_fu_10250_p2;
wire   [0:0] z0_113_fu_10232_p2;
wire   [0:0] z2_110_fu_10256_p2;
wire   [0:0] xor_ln45_290_fu_10262_p2;
wire   [0:0] xor_ln45_291_fu_10268_p2;
wire   [1:0] a1_330_fu_10178_p4;
wire   [1:0] b1_229_fu_10194_p4;
wire   [0:0] a0_324_fu_10282_p3;
wire   [1:0] a_390_fu_10290_p2;
wire   [0:0] b0_116_fu_10296_p3;
wire   [1:0] b_343_fu_10304_p2;
wire   [0:0] b0_115_fu_10324_p2;
wire   [0:0] a0_323_fu_10310_p2;
wire   [0:0] a1_332_fu_10316_p3;
wire   [0:0] b1_231_fu_10330_p3;
wire   [0:0] a_392_fu_10344_p2;
wire   [0:0] b_345_fu_10350_p2;
wire   [0:0] z1_113_fu_10356_p2;
wire   [0:0] z0_115_fu_10338_p2;
wire   [0:0] z2_111_fu_10362_p2;
wire   [0:0] xor_ln45_292_fu_10368_p2;
wire   [0:0] xor_ln45_293_fu_10374_p2;
wire   [0:0] a1_333_fu_10388_p3;
wire   [0:0] b1_232_fu_10396_p3;
wire   [0:0] a_396_fu_10410_p2;
wire   [0:0] b_349_fu_10416_p2;
wire   [0:0] z1_115_fu_10422_p2;
wire   [0:0] z0_116_fu_10404_p2;
wire   [0:0] z2_112_fu_10428_p2;
wire   [0:0] a1_191_fu_10434_p2;
wire   [0:0] a0_193_fu_10440_p2;
wire   [0:0] xor_ln28_47_fu_10454_p2;
wire   [1:0] z1_114_fu_10380_p3;
wire   [1:0] z0_114_fu_10274_p3;
wire   [1:0] z2_156_fu_10446_p3;
wire   [1:0] tmp_46_fu_10460_p3;
wire   [1:0] xor_ln45_297_fu_10474_p2;
wire   [1:0] xor_ln45_296_fu_10468_p2;
wire   [1:0] xor_ln45_298_fu_10480_p2;
wire   [1:0] xor_ln45_299_fu_10486_p2;
wire   [0:0] a1_335_fu_10520_p3;
wire   [0:0] b1_234_fu_10528_p3;
wire   [0:0] a_402_fu_10542_p2;
wire   [0:0] b_354_fu_10548_p2;
wire   [0:0] z1_117_fu_10554_p2;
wire   [0:0] z0_117_fu_10536_p2;
wire   [0:0] z2_114_fu_10560_p2;
wire   [0:0] xor_ln45_300_fu_10566_p2;
wire   [0:0] xor_ln45_301_fu_10572_p2;
wire   [1:0] a1_334_fu_10500_p4;
wire   [1:0] b1_233_fu_10510_p4;
wire   [0:0] a0_328_fu_10586_p3;
wire   [1:0] a_404_fu_10594_p2;
wire   [0:0] b0_120_fu_10600_p3;
wire   [1:0] b_356_fu_10608_p2;
wire   [0:0] b0_119_fu_10628_p2;
wire   [0:0] a0_327_fu_10614_p2;
wire   [0:0] a1_336_fu_10620_p3;
wire   [0:0] b1_235_fu_10634_p3;
wire   [0:0] a_406_fu_10648_p2;
wire   [0:0] b_358_fu_10654_p2;
wire   [0:0] z1_118_fu_10660_p2;
wire   [0:0] z0_119_fu_10642_p2;
wire   [0:0] z2_115_fu_10666_p2;
wire   [0:0] xor_ln45_302_fu_10672_p2;
wire   [0:0] xor_ln45_303_fu_10678_p2;
wire   [0:0] a1_337_fu_10692_p3;
wire   [0:0] b1_236_fu_10700_p3;
wire   [0:0] a_410_fu_10714_p2;
wire   [0:0] b_362_fu_10720_p2;
wire   [0:0] z1_120_fu_10726_p2;
wire   [0:0] z0_120_fu_10708_p2;
wire   [0:0] z2_116_fu_10732_p2;
wire   [0:0] a1_fu_10738_p2;
wire   [0:0] a0_198_fu_10744_p2;
wire   [0:0] xor_ln28_48_fu_10758_p2;
wire   [1:0] z1_119_fu_10684_p3;
wire   [1:0] z0_118_fu_10578_p3;
wire   [1:0] z2_157_fu_10750_p3;
wire   [1:0] tmp_47_fu_10764_p3;
wire   [1:0] xor_ln45_307_fu_10778_p2;
wire   [1:0] xor_ln45_306_fu_10772_p2;
wire   [1:0] a1_338_fu_10784_p2;
wire   [1:0] a0_199_fu_10790_p2;
wire   [0:0] a0_200_fu_10804_p1;
wire   [0:0] a1_197_fu_10808_p3;
wire   [0:0] xor_ln28_49_fu_10816_p2;
wire   [1:0] tmp_48_fu_10822_p3;
wire   [1:0] xor_ln28_50_fu_10830_p2;
wire   [3:0] z1_116_fu_10492_p3;
wire   [3:0] z0_112_fu_10116_p3;
wire   [3:0] z2_158_fu_10796_p3;
wire   [3:0] tmp_49_fu_10836_p3;
wire   [3:0] xor_ln45_311_fu_10850_p2;
wire   [3:0] xor_ln45_310_fu_10844_p2;
wire   [3:0] a1_339_fu_10856_p2;
wire   [3:0] a0_201_fu_10862_p2;
wire   [0:0] a0_203_fu_10890_p3;
wire   [0:0] a1_200_fu_10898_p3;
wire   [0:0] xor_ln28_51_fu_10906_p2;
wire   [1:0] a0_202_fu_10876_p1;
wire   [1:0] tmp_50_fu_10912_p3;
wire   [1:0] xor_ln28_52_fu_10920_p2;
wire   [1:0] a1_340_fu_10880_p4;
wire   [3:0] tmp_51_fu_10926_p3;
wire   [3:0] xor_ln28_53_fu_10934_p2;
wire   [7:0] z1_107_fu_9792_p3;
wire   [7:0] z0_94_fu_8580_p3;
wire   [7:0] z2_159_fu_10868_p3;
wire   [7:0] tmp_52_fu_10940_p3;
wire   [7:0] xor_ln45_315_fu_10954_p2;
wire   [7:0] xor_ln45_314_fu_10948_p2;
wire   [7:0] a1_341_fu_10960_p2;
wire   [7:0] a0_204_fu_10966_p2;
wire   [0:0] a0_207_fu_11014_p3;
wire   [0:0] a1_204_fu_11022_p3;
wire   [0:0] xor_ln28_54_fu_11030_p2;
wire   [1:0] a0_206_fu_10994_p4;
wire   [1:0] tmp_53_fu_11036_p3;
wire   [1:0] xor_ln28_55_fu_11044_p2;
wire   [1:0] a1_343_fu_11004_p4;
wire   [3:0] a0_205_fu_10980_p1;
wire   [3:0] tmp_54_fu_11050_p3;
wire   [3:0] xor_ln28_56_fu_11058_p2;
wire   [3:0] a1_342_fu_10984_p4;
wire   [7:0] tmp_55_fu_11064_p3;
wire   [7:0] xor_ln28_57_fu_11072_p2;
wire   [15:0] z1_80_fu_7484_p3;
wire   [15:0] z0_40_fu_3732_p3;
wire   [15:0] z2_160_fu_10972_p3;
wire   [15:0] tmp_56_fu_11078_p3;
wire   [15:0] xor_ln45_319_fu_11092_p2;
wire   [15:0] xor_ln45_318_fu_11086_p2;
wire   [15:0] xor_ln45_320_fu_11098_p2;
wire   [15:0] xor_ln45_321_fu_11104_p2;

assign a0_102_fu_4968_p2 = (z2_50_fu_4956_p2 ^ z0_53_fu_4932_p2);

assign a0_103_fu_5014_p2 = (z2_136_fu_4974_p3 ^ z0_51_fu_4802_p3);

assign a0_105_fu_5028_p1 = a1_265_fu_5008_p2[0:0];

assign a0_114_fu_5500_p2 = (z2_55_fu_5488_p2 ^ z0_58_fu_5464_p2);

assign a0_123_fu_5876_p2 = (z2_59_fu_5864_p2 ^ z0_63_fu_5840_p2);

assign a0_129_fu_6180_p2 = (z2_63_fu_6168_p2 ^ z0_67_fu_6144_p2);

assign a0_130_fu_6226_p2 = (z2_140_fu_6186_p3 ^ z0_65_fu_6014_p3);

assign a0_131_fu_6240_p1 = a1_279_fu_6220_p2[0:0];

assign a0_135_fu_6576_p2 = (z2_68_fu_6564_p2 ^ z0_71_fu_6540_p2);

assign a0_13_fu_912_p2 = (z2_6_fu_900_p2 ^ z0_8_fu_876_p2);

assign a0_140_fu_6952_p2 = (z2_72_fu_6940_p2 ^ z0_76_fu_6916_p2);

assign a0_144_fu_7256_p2 = (z2_76_fu_7244_p2 ^ z0_80_fu_7220_p2);

assign a0_145_fu_7302_p2 = (z2_144_fu_7262_p3 ^ z0_78_fu_7090_p3);

assign a0_146_fu_7316_p1 = a1_293_fu_7296_p2[0:0];

assign a0_147_fu_7374_p2 = (z2_145_fu_7308_p3 ^ z0_72_fu_6628_p3);

assign a0_148_fu_7388_p1 = a1_294_fu_7368_p2[1:0];

assign a0_149_fu_7402_p3 = a1_294_fu_7368_p2[32'd2];

assign a0_154_fu_7776_p2 = (z2_82_fu_7764_p2 ^ z0_84_fu_7740_p2);

assign a0_159_fu_8152_p2 = (z2_86_fu_8140_p2 ^ z0_89_fu_8116_p2);

assign a0_164_fu_8456_p2 = (z2_90_fu_8444_p2 ^ z0_93_fu_8420_p2);

assign a0_165_fu_8502_p2 = (z2_149_fu_8462_p3 ^ z0_91_fu_8290_p3);

assign a0_166_fu_8516_p1 = a1_310_fu_8496_p2[0:0];

assign a0_172_fu_8988_p2 = (z2_95_fu_8976_p2 ^ z0_98_fu_8952_p2);

assign a0_177_fu_9364_p2 = (z2_99_fu_9352_p2 ^ z0_103_fu_9328_p2);

assign a0_181_fu_9668_p2 = (z2_103_fu_9656_p2 ^ z0_107_fu_9632_p2);

assign a0_182_fu_9714_p2 = (z2_153_fu_9674_p3 ^ z0_105_fu_9502_p3);

assign a0_183_fu_9728_p1 = a1_324_fu_9708_p2[0:0];

assign a0_188_fu_10064_p2 = (z2_108_fu_10052_p2 ^ z0_111_fu_10028_p2);

assign a0_193_fu_10440_p2 = (z2_112_fu_10428_p2 ^ z0_116_fu_10404_p2);

assign a0_198_fu_10744_p2 = (z2_116_fu_10732_p2 ^ z0_120_fu_10708_p2);

assign a0_199_fu_10790_p2 = (z2_157_fu_10750_p3 ^ z0_118_fu_10578_p3);

assign a0_200_fu_10804_p1 = a1_338_fu_10784_p2[0:0];

assign a0_201_fu_10862_p2 = (z2_158_fu_10796_p3 ^ z0_112_fu_10116_p3);

assign a0_202_fu_10876_p1 = a1_339_fu_10856_p2[1:0];

assign a0_203_fu_10890_p3 = a1_339_fu_10856_p2[32'd2];

assign a0_204_fu_10966_p2 = (z2_159_fu_10868_p3 ^ z0_94_fu_8580_p3);

assign a0_205_fu_10980_p1 = a1_341_fu_10960_p2[3:0];

assign a0_206_fu_10994_p4 = {{a1_341_fu_10960_p2[5:4]}};

assign a0_207_fu_11014_p3 = a1_341_fu_10960_p2[32'd6];

assign a0_208_fu_160_p1 = a[15:0];

assign a0_209_fu_212_p1 = a[7:0];

assign a0_20_fu_1216_p2 = (z2_10_fu_1204_p2 ^ z0_12_fu_1180_p2);

assign a0_210_fu_248_p1 = a[3:0];

assign a0_211_fu_276_p1 = a[1:0];

assign a0_212_fu_304_p1 = a[0:0];

assign a0_213_fu_406_p2 = (a0_214_fu_378_p3 ^ a0_212_fu_304_p1);

assign a0_214_fu_378_p3 = a[32'd2];

assign a0_215_fu_644_p2 = (a0_219_fu_604_p4 ^ a0_211_fu_276_p1);

assign a0_216_fu_676_p2 = (a0_220_fu_596_p3 ^ a0_212_fu_304_p1);

assign a0_217_fu_782_p2 = (a0_218_fu_754_p3 ^ a0_216_fu_676_p2);

assign a0_218_fu_754_p3 = a_17_fu_614_p2[32'd2];

assign a0_219_fu_604_p4 = {{a[5:4]}};

assign a0_21_fu_1262_p2 = (z2_123_fu_1222_p3 ^ z0_10_fu_1050_p3);

assign a0_220_fu_596_p3 = a[32'd4];

assign a0_221_fu_1086_p2 = (a0_222_fu_1058_p3 ^ a0_220_fu_596_p3);

assign a0_222_fu_1058_p3 = a[32'd6];

assign a0_223_fu_1448_p2 = (a0_236_fu_1366_p4 ^ a0_210_fu_248_p1);

assign a0_224_fu_1480_p2 = (a0_237_fu_1356_p4 ^ a0_211_fu_276_p1);

assign a0_225_fu_1512_p2 = (a0_238_fu_1348_p3 ^ a0_212_fu_304_p1);

assign a0_226_fu_1618_p2 = (a0_227_fu_1590_p3 ^ a0_225_fu_1512_p2);

assign a0_227_fu_1590_p3 = a0_223_fu_1448_p2[32'd2];

assign a0_228_fu_1856_p2 = (a0_232_fu_1816_p4 ^ a0_224_fu_1480_p2);

assign a0_229_fu_1888_p2 = (a0_233_fu_1808_p3 ^ a0_225_fu_1512_p2);

assign a0_230_fu_1994_p2 = (a0_231_fu_1966_p3 ^ a0_229_fu_1888_p2);

assign a0_231_fu_1966_p3 = a_62_fu_1826_p2[32'd2];

assign a0_232_fu_1816_p4 = {{a_47_fu_1386_p2[5:4]}};

assign a0_233_fu_1808_p3 = a_47_fu_1386_p2[32'd4];

assign a0_234_fu_2298_p2 = (a0_235_fu_2270_p3 ^ a0_233_fu_1808_p3);

assign a0_235_fu_2270_p3 = a_47_fu_1386_p2[32'd6];

assign a0_236_fu_1366_p4 = {{a[11:8]}};

assign a0_237_fu_1356_p4 = {{a[9:8]}};

assign a0_238_fu_1348_p3 = a[32'd8];

assign a0_239_fu_2694_p2 = (a0_240_fu_2666_p3 ^ a0_238_fu_1348_p3);

assign a0_23_fu_1276_p1 = a1_220_fu_1256_p2[0:0];

assign a0_240_fu_2666_p3 = a[32'd10];

assign a0_241_fu_2932_p2 = (a0_245_fu_2892_p4 ^ a0_237_fu_1356_p4);

assign a0_242_fu_2964_p2 = (a0_246_fu_2884_p3 ^ a0_238_fu_1348_p3);

assign a0_243_fu_3070_p2 = (a0_244_fu_3042_p3 ^ a0_242_fu_2964_p2);

assign a0_244_fu_3042_p3 = a_107_fu_2902_p2[32'd2];

assign a0_245_fu_2892_p4 = {{a[13:12]}};

assign a0_246_fu_2884_p3 = a[32'd12];

assign a0_247_fu_3374_p2 = (a0_248_fu_3346_p3 ^ a0_246_fu_2884_p3);

assign a0_248_fu_3346_p3 = a[32'd14];

assign a0_249_fu_3934_p2 = (a0_289_fu_3768_p4 ^ a0_209_fu_212_p1);

assign a0_250_fu_3988_p2 = (a0_290_fu_3758_p4 ^ a0_210_fu_248_p1);

assign a0_251_fu_4020_p2 = (a0_291_fu_3748_p4 ^ a0_211_fu_276_p1);

assign a0_252_fu_4052_p2 = (a0_292_fu_3740_p3 ^ a0_212_fu_304_p1);

assign a0_253_fu_4158_p2 = (a0_254_fu_4130_p3 ^ a0_252_fu_4052_p2);

assign a0_254_fu_4130_p3 = a0_250_fu_3988_p2[32'd2];

assign a0_255_fu_4396_p2 = (a0_259_fu_4356_p4 ^ a0_251_fu_4020_p2);

assign a0_256_fu_4428_p2 = (a0_260_fu_4348_p3 ^ a0_252_fu_4052_p2);

assign a0_257_fu_4534_p2 = (a0_258_fu_4506_p3 ^ a0_256_fu_4428_p2);

assign a0_258_fu_4506_p3 = a_156_fu_4366_p2[32'd2];

assign a0_259_fu_4356_p4 = {{a0_249_fu_3934_p2[5:4]}};

assign a0_260_fu_4348_p3 = a0_249_fu_3934_p2[32'd4];

assign a0_261_fu_4838_p2 = (a0_262_fu_4810_p3 ^ a0_260_fu_4348_p3);

assign a0_262_fu_4810_p3 = a0_249_fu_3934_p2[32'd6];

assign a0_263_fu_5200_p2 = (a0_276_fu_5118_p4 ^ a0_250_fu_3988_p2);

assign a0_264_fu_5232_p2 = (a0_277_fu_5108_p4 ^ a0_251_fu_4020_p2);

assign a0_265_fu_5264_p2 = (a0_278_fu_5100_p3 ^ a0_252_fu_4052_p2);

assign a0_266_fu_5370_p2 = (a0_267_fu_5342_p3 ^ a0_265_fu_5264_p2);

assign a0_267_fu_5342_p3 = a0_263_fu_5200_p2[32'd2];

assign a0_268_fu_5608_p2 = (a0_272_fu_5568_p4 ^ a0_264_fu_5232_p2);

assign a0_269_fu_5640_p2 = (a0_273_fu_5560_p3 ^ a0_265_fu_5264_p2);

assign a0_270_fu_5746_p2 = (a0_271_fu_5718_p3 ^ a0_269_fu_5640_p2);

assign a0_271_fu_5718_p3 = a_201_fu_5578_p2[32'd2];

assign a0_272_fu_5568_p4 = {{a_186_fu_5138_p2[5:4]}};

assign a0_273_fu_5560_p3 = a_186_fu_5138_p2[32'd4];

assign a0_274_fu_6050_p2 = (a0_275_fu_6022_p3 ^ a0_273_fu_5560_p3);

assign a0_275_fu_6022_p3 = a_186_fu_5138_p2[32'd6];

assign a0_276_fu_5118_p4 = {{a_140_fu_3808_p2[11:8]}};

assign a0_277_fu_5108_p4 = {{a_140_fu_3808_p2[9:8]}};

assign a0_278_fu_5100_p3 = a_140_fu_3808_p2[32'd8];

assign a0_279_fu_6446_p2 = (a0_280_fu_6418_p3 ^ a0_278_fu_5100_p3);

assign a0_280_fu_6418_p3 = xor_ln43_44_fu_3826_p2[32'd10];

assign a0_281_fu_6684_p2 = (a0_285_fu_6644_p4 ^ a0_277_fu_5108_p4);

assign a0_282_fu_6716_p2 = (a0_286_fu_6636_p3 ^ a0_278_fu_5100_p3);

assign a0_283_fu_6822_p2 = (a0_284_fu_6794_p3 ^ a0_282_fu_6716_p2);

assign a0_284_fu_6794_p3 = a_246_fu_6654_p2[32'd2];

assign a0_285_fu_6644_p4 = {{a_140_fu_3808_p2[13:12]}};

assign a0_286_fu_6636_p3 = a_140_fu_3808_p2[32'd12];

assign a0_287_fu_7126_p2 = (a0_288_fu_7098_p3 ^ a0_286_fu_6636_p3);

assign a0_288_fu_7098_p3 = a_140_fu_3808_p2[32'd14];

assign a0_289_fu_3768_p4 = {{a[23:16]}};

assign a0_290_fu_3758_p4 = {{a[19:16]}};

assign a0_291_fu_3748_p4 = {{a[17:16]}};

assign a0_292_fu_3740_p3 = a[32'd16];

assign a0_293_fu_7646_p2 = (a0_294_fu_7618_p3 ^ a0_292_fu_3740_p3);

assign a0_294_fu_7618_p3 = a[32'd18];

assign a0_295_fu_7884_p2 = (a0_299_fu_7844_p4 ^ a0_291_fu_3748_p4);

assign a0_296_fu_7916_p2 = (a0_300_fu_7836_p3 ^ a0_292_fu_3740_p3);

assign a0_297_fu_8022_p2 = (a0_298_fu_7994_p3 ^ a0_296_fu_7916_p2);

assign a0_298_fu_7994_p3 = a_295_fu_7854_p2[32'd2];

assign a0_299_fu_7844_p4 = {{a[21:20]}};

assign a0_300_fu_7836_p3 = a[32'd20];

assign a0_301_fu_8326_p2 = (a0_302_fu_8298_p3 ^ a0_300_fu_7836_p3);

assign a0_302_fu_8298_p3 = a[32'd22];

assign a0_303_fu_8688_p2 = (a0_316_fu_8606_p4 ^ a0_290_fu_3758_p4);

assign a0_304_fu_8720_p2 = (a0_317_fu_8596_p4 ^ a0_291_fu_3748_p4);

assign a0_305_fu_8752_p2 = (a0_318_fu_8588_p3 ^ a0_292_fu_3740_p3);

assign a0_306_fu_8858_p2 = (a0_307_fu_8830_p3 ^ a0_305_fu_8752_p2);

assign a0_307_fu_8830_p3 = a0_303_fu_8688_p2[32'd2];

assign a0_308_fu_9096_p2 = (a0_312_fu_9056_p4 ^ a0_304_fu_8720_p2);

assign a0_309_fu_9128_p2 = (a0_313_fu_9048_p3 ^ a0_305_fu_8752_p2);

assign a0_310_fu_9234_p2 = (a0_311_fu_9206_p3 ^ a0_309_fu_9128_p2);

assign a0_311_fu_9206_p3 = a_340_fu_9066_p2[32'd2];

assign a0_312_fu_9056_p4 = {{a_325_fu_8626_p2[5:4]}};

assign a0_313_fu_9048_p3 = a_325_fu_8626_p2[32'd4];

assign a0_314_fu_9538_p2 = (a0_315_fu_9510_p3 ^ a0_313_fu_9048_p3);

assign a0_315_fu_9510_p3 = a_325_fu_8626_p2[32'd6];

assign a0_316_fu_8606_p4 = {{a[27:24]}};

assign a0_317_fu_8596_p4 = {{a[25:24]}};

assign a0_318_fu_8588_p3 = a[32'd24];

assign a0_319_fu_9934_p2 = (a0_320_fu_9906_p3 ^ a0_318_fu_8588_p3);

assign a0_320_fu_9906_p3 = a[32'd26];

assign a0_321_fu_10172_p2 = (a0_325_fu_10132_p4 ^ a0_317_fu_8596_p4);

assign a0_322_fu_10204_p2 = (a0_326_fu_10124_p3 ^ a0_318_fu_8588_p3);

assign a0_323_fu_10310_p2 = (a0_324_fu_10282_p3 ^ a0_322_fu_10204_p2);

assign a0_324_fu_10282_p3 = a_385_fu_10142_p2[32'd2];

assign a0_325_fu_10132_p4 = {{a[29:28]}};

assign a0_326_fu_10124_p3 = a[32'd28];

assign a0_327_fu_10614_p2 = (a0_328_fu_10586_p3 ^ a0_326_fu_10124_p3);

assign a0_328_fu_10586_p3 = a[32'd30];

assign a0_32_fu_1748_p2 = (z2_15_fu_1736_p2 ^ z0_17_fu_1712_p2);

assign a0_39_fu_2124_p2 = (z2_19_fu_2112_p2 ^ z0_22_fu_2088_p2);

assign a0_46_fu_2428_p2 = (z2_23_fu_2416_p2 ^ z0_26_fu_2392_p2);

assign a0_47_fu_2474_p2 = (z2_127_fu_2434_p3 ^ z0_24_fu_2262_p3);

assign a0_48_fu_2488_p1 = a1_234_fu_2468_p2[0:0];

assign a0_54_fu_2824_p2 = (z2_28_fu_2812_p2 ^ z0_30_fu_2788_p2);

assign a0_62_fu_3200_p2 = (z2_32_fu_3188_p2 ^ z0_35_fu_3164_p2);

assign a0_69_fu_3504_p2 = (z2_36_fu_3492_p2 ^ z0_39_fu_3468_p2);

assign a0_72_fu_3550_p2 = (z2_131_fu_3510_p3 ^ z0_37_fu_3338_p3);

assign a0_74_fu_3564_p1 = a1_248_fu_3544_p2[0:0];

assign a0_75_fu_3622_p2 = (z2_132_fu_3556_p3 ^ z0_31_fu_2876_p3);

assign a0_76_fu_3636_p1 = a1_249_fu_3616_p2[1:0];

assign a0_78_fu_3650_p3 = a1_249_fu_3616_p2[32'd2];

assign a0_90_fu_4288_p2 = (z2_42_fu_4276_p2 ^ z0_44_fu_4252_p2);

assign a0_97_fu_4664_p2 = (z2_46_fu_4652_p2 ^ z0_49_fu_4628_p2);

assign a0_fu_536_p2 = (z2_2_fu_524_p2 ^ z0_3_fu_500_p2);

assign a1_105_fu_5870_p2 = (z1_60_fu_5858_p2 ^ z0_63_fu_5840_p2);

assign a1_112_fu_6174_p2 = (z1_65_fu_6162_p2 ^ z0_67_fu_6144_p2);

assign a1_114_fu_6244_p3 = a1_279_fu_6220_p2[32'd1];

assign a1_120_fu_6570_p2 = (z1_70_fu_6558_p2 ^ z0_71_fu_6540_p2);

assign a1_126_fu_6946_p2 = (z1_74_fu_6934_p2 ^ z0_76_fu_6916_p2);

assign a1_133_fu_7250_p2 = (z1_79_fu_7238_p2 ^ z0_80_fu_7220_p2);

assign a1_135_fu_7320_p3 = a1_293_fu_7296_p2[32'd1];

assign a1_138_fu_7410_p3 = a1_294_fu_7368_p2[32'd3];

assign a1_147_fu_7770_p2 = (z1_84_fu_7758_p2 ^ z0_84_fu_7740_p2);

assign a1_153_fu_8146_p2 = (z1_88_fu_8134_p2 ^ z0_89_fu_8116_p2);

assign a1_159_fu_8450_p2 = (z1_93_fu_8438_p2 ^ z0_93_fu_8420_p2);

assign a1_15_fu_906_p2 = (z1_7_fu_894_p2 ^ z0_8_fu_876_p2);

assign a1_161_fu_8520_p3 = a1_310_fu_8496_p2[32'd1];

assign a1_168_fu_8982_p2 = (z1_97_fu_8970_p2 ^ z0_98_fu_8952_p2);

assign a1_173_fu_9358_p2 = (z1_101_fu_9346_p2 ^ z0_103_fu_9328_p2);

assign a1_178_fu_9662_p2 = (z1_106_fu_9650_p2 ^ z0_107_fu_9632_p2);

assign a1_180_fu_9732_p3 = a1_324_fu_9708_p2[32'd1];

assign a1_186_fu_10058_p2 = (z1_111_fu_10046_p2 ^ z0_111_fu_10028_p2);

assign a1_191_fu_10434_p2 = (z1_115_fu_10422_p2 ^ z0_116_fu_10404_p2);

assign a1_197_fu_10808_p3 = a1_338_fu_10784_p2[32'd1];

assign a1_200_fu_10898_p3 = a1_339_fu_10856_p2[32'd3];

assign a1_204_fu_11022_p3 = a1_341_fu_10960_p2[32'd7];

assign a1_205_fu_176_p4 = {{a[31:16]}};

assign a1_206_fu_220_p4 = {{a[15:8]}};

assign a1_207_fu_252_p4 = {{a[7:4]}};

assign a1_208_fu_280_p4 = {{a[3:2]}};

assign a1_209_fu_308_p3 = a[32'd1];

assign a1_210_fu_412_p3 = a_8_fu_386_p2[32'd1];

assign a1_211_fu_484_p3 = a[32'd3];

assign a1_212_fu_650_p4 = {{a_17_fu_614_p2[3:2]}};

assign a1_213_fu_682_p3 = a0_215_fu_644_p2[32'd1];

assign a1_214_fu_788_p3 = a_22_fu_762_p2[32'd1];

assign a1_215_fu_860_p3 = a_17_fu_614_p2[32'd3];

assign a1_216_fu_972_p4 = {{a[7:6]}};

assign a1_217_fu_992_p3 = a[32'd5];

assign a1_218_fu_1092_p3 = a_36_fu_1066_p2[32'd1];

assign a1_219_fu_1164_p3 = a[32'd7];

assign a1_21_fu_1210_p2 = (z1_12_fu_1198_p2 ^ z0_12_fu_1180_p2);

assign a1_220_fu_1256_p2 = (xor_ln45_27_fu_1250_p2 ^ xor_ln45_26_fu_1244_p2);

assign a1_221_fu_1454_p4 = {{a_47_fu_1386_p2[7:4]}};

assign a1_222_fu_1486_p4 = {{a0_223_fu_1448_p2[3:2]}};

assign a1_223_fu_1518_p3 = a0_224_fu_1480_p2[32'd1];

assign a1_224_fu_1624_p3 = a_53_fu_1598_p2[32'd1];

assign a1_225_fu_1696_p3 = a0_223_fu_1448_p2[32'd3];

assign a1_226_fu_1862_p4 = {{a_62_fu_1826_p2[3:2]}};

assign a1_227_fu_1894_p3 = a0_228_fu_1856_p2[32'd1];

assign a1_228_fu_2000_p3 = a_67_fu_1974_p2[32'd1];

assign a1_229_fu_2072_p3 = a_62_fu_1826_p2[32'd3];

assign a1_230_fu_2184_p4 = {{a_47_fu_1386_p2[7:6]}};

assign a1_231_fu_2204_p3 = xor_ln43_14_fu_1392_p2[32'd5];

assign a1_232_fu_2304_p3 = a_81_fu_2278_p2[32'd1];

assign a1_233_fu_2376_p3 = a_47_fu_1386_p2[32'd7];

assign a1_234_fu_2468_p2 = (xor_ln45_61_fu_2462_p2 ^ xor_ln45_60_fu_2456_p2);

assign a1_235_fu_2560_p4 = {{a[15:12]}};

assign a1_236_fu_2580_p4 = {{a[11:10]}};

assign a1_237_fu_2600_p3 = a[32'd9];

assign a1_238_fu_2700_p3 = a_98_fu_2674_p2[32'd1];

assign a1_239_fu_2772_p3 = a[32'd11];

assign a1_23_fu_1280_p3 = a1_220_fu_1256_p2[32'd1];

assign a1_240_fu_2938_p4 = {{a_107_fu_2902_p2[3:2]}};

assign a1_241_fu_2970_p3 = a0_241_fu_2932_p2[32'd1];

assign a1_242_fu_3076_p3 = a_112_fu_3050_p2[32'd1];

assign a1_243_fu_3148_p3 = a_107_fu_2902_p2[32'd3];

assign a1_244_fu_3260_p4 = {{a[15:14]}};

assign a1_245_fu_3280_p3 = a[32'd13];

assign a1_246_fu_3380_p3 = a_126_fu_3354_p2[32'd1];

assign a1_247_fu_3452_p3 = a[32'd15];

assign a1_248_fu_3544_p2 = (xor_ln45_95_fu_3538_p2 ^ xor_ln45_94_fu_3532_p2);

assign a1_249_fu_3616_p2 = (xor_ln45_99_fu_3610_p2 ^ xor_ln45_98_fu_3604_p2);

assign a1_250_fu_3640_p4 = {{a1_249_fu_3616_p2[3:2]}};

assign a1_251_fu_3946_p4 = {{a_140_fu_3808_p2[15:8]}};

assign a1_252_fu_3994_p4 = {{a0_249_fu_3934_p2[7:4]}};

assign a1_253_fu_4026_p4 = {{a0_250_fu_3988_p2[3:2]}};

assign a1_254_fu_4058_p3 = a0_251_fu_4020_p2[32'd1];

assign a1_255_fu_4164_p3 = a_147_fu_4138_p2[32'd1];

assign a1_256_fu_4236_p3 = a0_250_fu_3988_p2[32'd3];

assign a1_257_fu_4402_p4 = {{a_156_fu_4366_p2[3:2]}};

assign a1_258_fu_4434_p3 = a0_255_fu_4396_p2[32'd1];

assign a1_259_fu_4540_p3 = a_161_fu_4514_p2[32'd1];

assign a1_260_fu_4612_p3 = a_156_fu_4366_p2[32'd3];

assign a1_261_fu_4724_p4 = {{a0_249_fu_3934_p2[7:6]}};

assign a1_262_fu_4744_p3 = xor_ln38_1_fu_3940_p2[32'd5];

assign a1_263_fu_4844_p3 = a_175_fu_4818_p2[32'd1];

assign a1_264_fu_4916_p3 = a0_249_fu_3934_p2[32'd7];

assign a1_265_fu_5008_p2 = (xor_ln45_133_fu_5002_p2 ^ xor_ln45_132_fu_4996_p2);

assign a1_266_fu_5206_p4 = {{a_186_fu_5138_p2[7:4]}};

assign a1_267_fu_5238_p4 = {{a0_263_fu_5200_p2[3:2]}};

assign a1_268_fu_5270_p3 = a0_264_fu_5232_p2[32'd1];

assign a1_269_fu_5376_p3 = a_192_fu_5350_p2[32'd1];

assign a1_270_fu_5448_p3 = a0_263_fu_5200_p2[32'd3];

assign a1_271_fu_5614_p4 = {{a_201_fu_5578_p2[3:2]}};

assign a1_272_fu_5646_p3 = a0_268_fu_5608_p2[32'd1];

assign a1_273_fu_5752_p3 = a_206_fu_5726_p2[32'd1];

assign a1_274_fu_5824_p3 = a_201_fu_5578_p2[32'd3];

assign a1_275_fu_5936_p4 = {{a_186_fu_5138_p2[7:6]}};

assign a1_276_fu_5956_p3 = xor_ln43_59_fu_5144_p2[32'd5];

assign a1_277_fu_6056_p3 = a_220_fu_6030_p2[32'd1];

assign a1_278_fu_6128_p3 = a_186_fu_5138_p2[32'd7];

assign a1_279_fu_6220_p2 = (xor_ln45_167_fu_6214_p2 ^ xor_ln45_166_fu_6208_p2);

assign a1_280_fu_6312_p4 = {{a_140_fu_3808_p2[15:12]}};

assign a1_281_fu_6332_p4 = {{xor_ln43_44_fu_3826_p2[11:10]}};

assign a1_282_fu_6352_p3 = xor_ln43_43_fu_3820_p2[32'd9];

assign a1_283_fu_6452_p3 = a_237_fu_6426_p2[32'd1];

assign a1_284_fu_6524_p3 = xor_ln43_44_fu_3826_p2[32'd11];

assign a1_285_fu_6690_p4 = {{a_246_fu_6654_p2[3:2]}};

assign a1_286_fu_6722_p3 = a0_281_fu_6684_p2[32'd1];

assign a1_287_fu_6828_p3 = a_251_fu_6802_p2[32'd1];

assign a1_288_fu_6900_p3 = a_246_fu_6654_p2[32'd3];

assign a1_289_fu_7012_p4 = {{a_140_fu_3808_p2[15:14]}};

assign a1_290_fu_7032_p3 = xor_ln43_42_fu_3814_p2[32'd13];

assign a1_291_fu_7132_p3 = a_265_fu_7106_p2[32'd1];

assign a1_292_fu_7204_p3 = a_140_fu_3808_p2[32'd15];

assign a1_293_fu_7296_p2 = (xor_ln45_201_fu_7290_p2 ^ xor_ln45_200_fu_7284_p2);

assign a1_294_fu_7368_p2 = (xor_ln45_205_fu_7362_p2 ^ xor_ln45_204_fu_7356_p2);

assign a1_295_fu_7392_p4 = {{a1_294_fu_7368_p2[3:2]}};

assign a1_296_fu_7492_p4 = {{a[31:24]}};

assign a1_297_fu_7512_p4 = {{a[23:20]}};

assign a1_298_fu_7532_p4 = {{a[19:18]}};

assign a1_299_fu_7552_p3 = a[32'd17];

assign a1_300_fu_7652_p3 = a_286_fu_7626_p2[32'd1];

assign a1_301_fu_7724_p3 = a[32'd19];

assign a1_302_fu_7890_p4 = {{a_295_fu_7854_p2[3:2]}};

assign a1_303_fu_7922_p3 = a0_295_fu_7884_p2[32'd1];

assign a1_304_fu_8028_p3 = a_300_fu_8002_p2[32'd1];

assign a1_305_fu_8100_p3 = a_295_fu_7854_p2[32'd3];

assign a1_306_fu_8212_p4 = {{a[23:22]}};

assign a1_307_fu_8232_p3 = a[32'd21];

assign a1_308_fu_8332_p3 = a_314_fu_8306_p2[32'd1];

assign a1_309_fu_8404_p3 = a[32'd23];

assign a1_310_fu_8496_p2 = (xor_ln45_239_fu_8490_p2 ^ xor_ln45_238_fu_8484_p2);

assign a1_311_fu_8694_p4 = {{a_325_fu_8626_p2[7:4]}};

assign a1_312_fu_8726_p4 = {{a0_303_fu_8688_p2[3:2]}};

assign a1_313_fu_8758_p3 = a0_304_fu_8720_p2[32'd1];

assign a1_314_fu_8864_p3 = a_331_fu_8838_p2[32'd1];

assign a1_315_fu_8936_p3 = a0_303_fu_8688_p2[32'd3];

assign a1_316_fu_9102_p4 = {{a_340_fu_9066_p2[3:2]}};

assign a1_317_fu_9134_p3 = a0_308_fu_9096_p2[32'd1];

assign a1_318_fu_9240_p3 = a_345_fu_9214_p2[32'd1];

assign a1_319_fu_9312_p3 = a_340_fu_9066_p2[32'd3];

assign a1_31_fu_1742_p2 = (z1_16_fu_1730_p2 ^ z0_17_fu_1712_p2);

assign a1_320_fu_9424_p4 = {{a_325_fu_8626_p2[7:6]}};

assign a1_321_fu_9444_p3 = xor_ln43_100_fu_8632_p2[32'd5];

assign a1_322_fu_9544_p3 = a_359_fu_9518_p2[32'd1];

assign a1_323_fu_9616_p3 = a_325_fu_8626_p2[32'd7];

assign a1_324_fu_9708_p2 = (xor_ln45_273_fu_9702_p2 ^ xor_ln45_272_fu_9696_p2);

assign a1_325_fu_9800_p4 = {{a[31:28]}};

assign a1_326_fu_9820_p4 = {{a[27:26]}};

assign a1_327_fu_9840_p3 = a[32'd25];

assign a1_328_fu_9940_p3 = a_376_fu_9914_p2[32'd1];

assign a1_329_fu_10012_p3 = a[32'd27];

assign a1_330_fu_10178_p4 = {{a_385_fu_10142_p2[3:2]}};

assign a1_331_fu_10210_p3 = a0_321_fu_10172_p2[32'd1];

assign a1_332_fu_10316_p3 = a_390_fu_10290_p2[32'd1];

assign a1_333_fu_10388_p3 = a_385_fu_10142_p2[32'd3];

assign a1_334_fu_10500_p4 = {{a[31:30]}};

assign a1_335_fu_10520_p3 = a[32'd29];

assign a1_336_fu_10620_p3 = a_404_fu_10594_p2[32'd1];

assign a1_337_fu_10692_p3 = a[32'd31];

assign a1_338_fu_10784_p2 = (xor_ln45_307_fu_10778_p2 ^ xor_ln45_306_fu_10772_p2);

assign a1_339_fu_10856_p2 = (xor_ln45_311_fu_10850_p2 ^ xor_ln45_310_fu_10844_p2);

assign a1_340_fu_10880_p4 = {{a1_339_fu_10856_p2[3:2]}};

assign a1_341_fu_10960_p2 = (xor_ln45_315_fu_10954_p2 ^ xor_ln45_314_fu_10948_p2);

assign a1_342_fu_10984_p4 = {{a1_341_fu_10960_p2[7:4]}};

assign a1_343_fu_11004_p4 = {{a1_341_fu_10960_p2[7:6]}};

assign a1_37_fu_2118_p2 = (z1_20_fu_2106_p2 ^ z0_22_fu_2088_p2);

assign a1_42_fu_2422_p2 = (z1_25_fu_2410_p2 ^ z0_26_fu_2392_p2);

assign a1_45_fu_2492_p3 = a1_234_fu_2468_p2[32'd1];

assign a1_52_fu_2818_p2 = (z1_30_fu_2806_p2 ^ z0_30_fu_2788_p2);

assign a1_58_fu_3194_p2 = (z1_34_fu_3182_p2 ^ z0_35_fu_3164_p2);

assign a1_63_fu_3498_p2 = (z1_39_fu_3486_p2 ^ z0_39_fu_3468_p2);

assign a1_66_fu_3568_p3 = a1_248_fu_3544_p2[32'd1];

assign a1_69_fu_3658_p3 = a1_249_fu_3616_p2[32'd3];

assign a1_78_fu_4282_p2 = (z1_43_fu_4270_p2 ^ z0_44_fu_4252_p2);

assign a1_84_fu_4658_p2 = (z1_47_fu_4646_p2 ^ z0_49_fu_4628_p2);

assign a1_90_fu_4962_p2 = (z1_52_fu_4950_p2 ^ z0_53_fu_4932_p2);

assign a1_92_fu_5032_p3 = a1_265_fu_5008_p2[32'd1];

assign a1_99_fu_5494_p2 = (z1_56_fu_5482_p2 ^ z0_58_fu_5464_p2);

assign a1_9_fu_530_p2 = (z1_3_fu_518_p2 ^ z0_3_fu_500_p2);

assign a1_fu_10738_p2 = (z1_120_fu_10726_p2 ^ z0_120_fu_10708_p2);

assign a_100_fu_2728_p2 = (a1_238_fu_2700_p3 ^ a0_239_fu_2694_p2);

assign a_104_fu_2794_p2 = (a1_239_fu_2772_p3 ^ a0_240_fu_2666_p3);

assign a_107_fu_2902_p2 = (a1_235_fu_2560_p4 ^ a0_236_fu_1366_p4);

assign a_10_fu_440_p2 = (a1_210_fu_412_p3 ^ a0_213_fu_406_p2);

assign a_110_fu_2998_p2 = (a1_241_fu_2970_p3 ^ a0_242_fu_2964_p2);

assign a_112_fu_3050_p2 = (a1_240_fu_2938_p4 ^ a0_241_fu_2932_p2);

assign a_114_fu_3104_p2 = (a1_242_fu_3076_p3 ^ a0_243_fu_3070_p2);

assign a_118_fu_3170_p2 = (a1_243_fu_3148_p3 ^ a0_244_fu_3042_p3);

assign a_124_fu_3302_p2 = (a1_245_fu_3280_p3 ^ a0_246_fu_2884_p3);

assign a_126_fu_3354_p2 = (a1_244_fu_3260_p4 ^ a0_245_fu_2892_p4);

assign a_128_fu_3408_p2 = (a1_246_fu_3380_p3 ^ a0_247_fu_3374_p2);

assign a_132_fu_3474_p2 = (a1_247_fu_3452_p3 ^ a0_248_fu_3346_p3);

assign a_140_fu_3808_p2 = (a1_205_fu_176_p4 ^ a0_208_fu_160_p1);

assign a_145_fu_4086_p2 = (a1_254_fu_4058_p3 ^ a0_252_fu_4052_p2);

assign a_147_fu_4138_p2 = (a1_253_fu_4026_p4 ^ a0_251_fu_4020_p2);

assign a_149_fu_4192_p2 = (a1_255_fu_4164_p3 ^ a0_253_fu_4158_p2);

assign a_14_fu_506_p2 = (a1_211_fu_484_p3 ^ a0_214_fu_378_p3);

assign a_153_fu_4258_p2 = (a1_256_fu_4236_p3 ^ a0_254_fu_4130_p3);

assign a_156_fu_4366_p2 = (a1_252_fu_3994_p4 ^ a0_250_fu_3988_p2);

assign a_159_fu_4462_p2 = (a1_258_fu_4434_p3 ^ a0_256_fu_4428_p2);

assign a_161_fu_4514_p2 = (a1_257_fu_4402_p4 ^ a0_255_fu_4396_p2);

assign a_163_fu_4568_p2 = (a1_259_fu_4540_p3 ^ a0_257_fu_4534_p2);

assign a_167_fu_4634_p2 = (a1_260_fu_4612_p3 ^ a0_258_fu_4506_p3);

assign a_173_fu_4766_p2 = (a1_262_fu_4744_p3 ^ a0_260_fu_4348_p3);

assign a_175_fu_4818_p2 = (a1_261_fu_4724_p4 ^ a0_259_fu_4356_p4);

assign a_177_fu_4872_p2 = (a1_263_fu_4844_p3 ^ a0_261_fu_4838_p2);

assign a_17_fu_614_p2 = (a1_207_fu_252_p4 ^ a0_210_fu_248_p1);

assign a_181_fu_4938_p2 = (a1_264_fu_4916_p3 ^ a0_262_fu_4810_p3);

assign a_186_fu_5138_p2 = (a1_251_fu_3946_p4 ^ a0_249_fu_3934_p2);

assign a_190_fu_5298_p2 = (a1_268_fu_5270_p3 ^ a0_265_fu_5264_p2);

assign a_192_fu_5350_p2 = (a1_267_fu_5238_p4 ^ a0_264_fu_5232_p2);

assign a_194_fu_5404_p2 = (a1_269_fu_5376_p3 ^ a0_266_fu_5370_p2);

assign a_198_fu_5470_p2 = (a1_270_fu_5448_p3 ^ a0_267_fu_5342_p3);

assign a_201_fu_5578_p2 = (a1_266_fu_5206_p4 ^ a0_263_fu_5200_p2);

assign a_204_fu_5674_p2 = (a1_272_fu_5646_p3 ^ a0_269_fu_5640_p2);

assign a_206_fu_5726_p2 = (a1_271_fu_5614_p4 ^ a0_268_fu_5608_p2);

assign a_208_fu_5780_p2 = (a1_273_fu_5752_p3 ^ a0_270_fu_5746_p2);

assign a_20_fu_710_p2 = (a1_213_fu_682_p3 ^ a0_216_fu_676_p2);

assign a_212_fu_5846_p2 = (a1_274_fu_5824_p3 ^ a0_271_fu_5718_p3);

assign a_218_fu_5978_p2 = (a1_276_fu_5956_p3 ^ a0_273_fu_5560_p3);

assign a_220_fu_6030_p2 = (a1_275_fu_5936_p4 ^ a0_272_fu_5568_p4);

assign a_222_fu_6084_p2 = (a1_277_fu_6056_p3 ^ a0_274_fu_6050_p2);

assign a_226_fu_6150_p2 = (a1_278_fu_6128_p3 ^ a0_275_fu_6022_p3);

assign a_22_fu_762_p2 = (a1_212_fu_650_p4 ^ a0_215_fu_644_p2);

assign a_235_fu_6374_p2 = (a1_282_fu_6352_p3 ^ a0_278_fu_5100_p3);

assign a_237_fu_6426_p2 = (a1_281_fu_6332_p4 ^ a0_277_fu_5108_p4);

assign a_239_fu_6480_p2 = (a1_283_fu_6452_p3 ^ a0_279_fu_6446_p2);

assign a_243_fu_6546_p2 = (a1_284_fu_6524_p3 ^ a0_280_fu_6418_p3);

assign a_246_fu_6654_p2 = (a1_280_fu_6312_p4 ^ a0_276_fu_5118_p4);

assign a_249_fu_6750_p2 = (a1_286_fu_6722_p3 ^ a0_282_fu_6716_p2);

assign a_24_fu_816_p2 = (a1_214_fu_788_p3 ^ a0_217_fu_782_p2);

assign a_251_fu_6802_p2 = (a1_285_fu_6690_p4 ^ a0_281_fu_6684_p2);

assign a_253_fu_6856_p2 = (a1_287_fu_6828_p3 ^ a0_283_fu_6822_p2);

assign a_257_fu_6922_p2 = (a1_288_fu_6900_p3 ^ a0_284_fu_6794_p3);

assign a_263_fu_7054_p2 = (a1_290_fu_7032_p3 ^ a0_286_fu_6636_p3);

assign a_265_fu_7106_p2 = (a1_289_fu_7012_p4 ^ a0_285_fu_6644_p4);

assign a_267_fu_7160_p2 = (a1_291_fu_7132_p3 ^ a0_287_fu_7126_p2);

assign a_271_fu_7226_p2 = (a1_292_fu_7204_p3 ^ a0_288_fu_7098_p3);

assign a_284_fu_7574_p2 = (a1_299_fu_7552_p3 ^ a0_292_fu_3740_p3);

assign a_286_fu_7626_p2 = (a1_298_fu_7532_p4 ^ a0_291_fu_3748_p4);

assign a_288_fu_7680_p2 = (a1_300_fu_7652_p3 ^ a0_293_fu_7646_p2);

assign a_28_fu_882_p2 = (a1_215_fu_860_p3 ^ a0_218_fu_754_p3);

assign a_292_fu_7746_p2 = (a1_301_fu_7724_p3 ^ a0_294_fu_7618_p3);

assign a_295_fu_7854_p2 = (a1_297_fu_7512_p4 ^ a0_290_fu_3758_p4);

assign a_298_fu_7950_p2 = (a1_303_fu_7922_p3 ^ a0_296_fu_7916_p2);

assign a_300_fu_8002_p2 = (a1_302_fu_7890_p4 ^ a0_295_fu_7884_p2);

assign a_302_fu_8056_p2 = (a1_304_fu_8028_p3 ^ a0_297_fu_8022_p2);

assign a_306_fu_8122_p2 = (a1_305_fu_8100_p3 ^ a0_298_fu_7994_p3);

assign a_312_fu_8254_p2 = (a1_307_fu_8232_p3 ^ a0_300_fu_7836_p3);

assign a_314_fu_8306_p2 = (a1_306_fu_8212_p4 ^ a0_299_fu_7844_p4);

assign a_316_fu_8360_p2 = (a1_308_fu_8332_p3 ^ a0_301_fu_8326_p2);

assign a_320_fu_8426_p2 = (a1_309_fu_8404_p3 ^ a0_302_fu_8298_p3);

assign a_325_fu_8626_p2 = (a1_296_fu_7492_p4 ^ a0_289_fu_3768_p4);

assign a_329_fu_8786_p2 = (a1_313_fu_8758_p3 ^ a0_305_fu_8752_p2);

assign a_331_fu_8838_p2 = (a1_312_fu_8726_p4 ^ a0_304_fu_8720_p2);

assign a_333_fu_8892_p2 = (a1_314_fu_8864_p3 ^ a0_306_fu_8858_p2);

assign a_337_fu_8958_p2 = (a1_315_fu_8936_p3 ^ a0_307_fu_8830_p3);

assign a_340_fu_9066_p2 = (a1_311_fu_8694_p4 ^ a0_303_fu_8688_p2);

assign a_343_fu_9162_p2 = (a1_317_fu_9134_p3 ^ a0_309_fu_9128_p2);

assign a_345_fu_9214_p2 = (a1_316_fu_9102_p4 ^ a0_308_fu_9096_p2);

assign a_347_fu_9268_p2 = (a1_318_fu_9240_p3 ^ a0_310_fu_9234_p2);

assign a_34_fu_1014_p2 = (a1_217_fu_992_p3 ^ a0_220_fu_596_p3);

assign a_351_fu_9334_p2 = (a1_319_fu_9312_p3 ^ a0_311_fu_9206_p3);

assign a_357_fu_9466_p2 = (a1_321_fu_9444_p3 ^ a0_313_fu_9048_p3);

assign a_359_fu_9518_p2 = (a1_320_fu_9424_p4 ^ a0_312_fu_9056_p4);

assign a_361_fu_9572_p2 = (a1_322_fu_9544_p3 ^ a0_314_fu_9538_p2);

assign a_365_fu_9638_p2 = (a1_323_fu_9616_p3 ^ a0_315_fu_9510_p3);

assign a_36_fu_1066_p2 = (a1_216_fu_972_p4 ^ a0_219_fu_604_p4);

assign a_374_fu_9862_p2 = (a1_327_fu_9840_p3 ^ a0_318_fu_8588_p3);

assign a_376_fu_9914_p2 = (a1_326_fu_9820_p4 ^ a0_317_fu_8596_p4);

assign a_378_fu_9968_p2 = (a1_328_fu_9940_p3 ^ a0_319_fu_9934_p2);

assign a_382_fu_10034_p2 = (a1_329_fu_10012_p3 ^ a0_320_fu_9906_p3);

assign a_385_fu_10142_p2 = (a1_325_fu_9800_p4 ^ a0_316_fu_8606_p4);

assign a_388_fu_10238_p2 = (a1_331_fu_10210_p3 ^ a0_322_fu_10204_p2);

assign a_38_fu_1120_p2 = (a1_218_fu_1092_p3 ^ a0_221_fu_1086_p2);

assign a_390_fu_10290_p2 = (a1_330_fu_10178_p4 ^ a0_321_fu_10172_p2);

assign a_392_fu_10344_p2 = (a1_332_fu_10316_p3 ^ a0_323_fu_10310_p2);

assign a_396_fu_10410_p2 = (a1_333_fu_10388_p3 ^ a0_324_fu_10282_p3);

assign a_402_fu_10542_p2 = (a1_335_fu_10520_p3 ^ a0_326_fu_10124_p3);

assign a_404_fu_10594_p2 = (a1_334_fu_10500_p4 ^ a0_325_fu_10132_p4);

assign a_406_fu_10648_p2 = (a1_336_fu_10620_p3 ^ a0_327_fu_10614_p2);

assign a_410_fu_10714_p2 = (a1_337_fu_10692_p3 ^ a0_328_fu_10586_p3);

assign a_42_fu_1186_p2 = (a1_219_fu_1164_p3 ^ a0_222_fu_1058_p3);

assign a_47_fu_1386_p2 = (a1_206_fu_220_p4 ^ a0_209_fu_212_p1);

assign a_51_fu_1546_p2 = (a1_223_fu_1518_p3 ^ a0_225_fu_1512_p2);

assign a_53_fu_1598_p2 = (a1_222_fu_1486_p4 ^ a0_224_fu_1480_p2);

assign a_55_fu_1652_p2 = (a1_224_fu_1624_p3 ^ a0_226_fu_1618_p2);

assign a_59_fu_1718_p2 = (a1_225_fu_1696_p3 ^ a0_227_fu_1590_p3);

assign a_62_fu_1826_p2 = (a1_221_fu_1454_p4 ^ a0_223_fu_1448_p2);

assign a_65_fu_1922_p2 = (a1_227_fu_1894_p3 ^ a0_229_fu_1888_p2);

assign a_67_fu_1974_p2 = (a1_226_fu_1862_p4 ^ a0_228_fu_1856_p2);

assign a_69_fu_2028_p2 = (a1_228_fu_2000_p3 ^ a0_230_fu_1994_p2);

assign a_6_fu_334_p2 = (a1_209_fu_308_p3 ^ a0_212_fu_304_p1);

assign a_73_fu_2094_p2 = (a1_229_fu_2072_p3 ^ a0_231_fu_1966_p3);

assign a_79_fu_2226_p2 = (a1_231_fu_2204_p3 ^ a0_233_fu_1808_p3);

assign a_81_fu_2278_p2 = (a1_230_fu_2184_p4 ^ a0_232_fu_1816_p4);

assign a_83_fu_2332_p2 = (a1_232_fu_2304_p3 ^ a0_234_fu_2298_p2);

assign a_87_fu_2398_p2 = (a1_233_fu_2376_p3 ^ a0_235_fu_2270_p3);

assign a_8_fu_386_p2 = (a1_208_fu_280_p4 ^ a0_211_fu_276_p1);

assign a_96_fu_2622_p2 = (a1_237_fu_2600_p3 ^ a0_238_fu_1348_p3);

assign a_98_fu_2674_p2 = (a1_236_fu_2580_p4 ^ a0_237_fu_1356_p4);

assign b0_100_fu_9112_p2 = (b0_96_fu_8736_p2 ^ b0_104_fu_9080_p4);

assign b0_101_fu_9142_p2 = (b0_97_fu_8766_p2 ^ b0_105_fu_9072_p3);

assign b0_102_fu_9248_p2 = (b0_103_fu_9220_p3 ^ b0_101_fu_9142_p2);

assign b0_103_fu_9220_p3 = b_298_fu_9090_p2[32'd2];

assign b0_104_fu_9080_p4 = {{b_284_fu_8676_p2[5:4]}};

assign b0_105_fu_9072_p3 = b_284_fu_8676_p2[32'd4];

assign b0_106_fu_9552_p2 = (b0_107_fu_9524_p3 ^ b0_105_fu_9072_p3);

assign b0_107_fu_9524_p3 = b_284_fu_8676_p2[32'd6];

assign b0_108_fu_8656_p4 = {{b[27:24]}};

assign b0_109_fu_8646_p4 = {{b[25:24]}};

assign b0_10_fu_768_p3 = b_16_fu_638_p2[32'd2];

assign b0_110_fu_8638_p3 = b[32'd24];

assign b0_111_fu_9948_p2 = (b0_112_fu_9920_p3 ^ b0_110_fu_8638_p3);

assign b0_112_fu_9920_p3 = b[32'd26];

assign b0_113_fu_10188_p2 = (b0_117_fu_10156_p4 ^ b0_109_fu_8646_p4);

assign b0_114_fu_10218_p2 = (b0_118_fu_10148_p3 ^ b0_110_fu_8638_p3);

assign b0_115_fu_10324_p2 = (b0_116_fu_10296_p3 ^ b0_114_fu_10218_p2);

assign b0_116_fu_10296_p3 = b_338_fu_10166_p2[32'd2];

assign b0_117_fu_10156_p4 = {{b[29:28]}};

assign b0_118_fu_10148_p3 = b[32'd28];

assign b0_119_fu_10628_p2 = (b0_120_fu_10600_p3 ^ b0_118_fu_10148_p3);

assign b0_11_fu_628_p4 = {{b[5:4]}};

assign b0_120_fu_10600_p3 = b[32'd30];

assign b0_12_fu_620_p3 = b[32'd4];

assign b0_13_fu_1100_p2 = (b0_14_fu_1072_p3 ^ b0_12_fu_620_p3);

assign b0_14_fu_1072_p3 = b[32'd6];

assign b0_15_fu_1464_p2 = (b0_2_fu_262_p1 ^ b0_28_fu_1416_p4);

assign b0_16_fu_1496_p2 = (b0_3_fu_290_p1 ^ b0_29_fu_1406_p4);

assign b0_17_fu_1526_p2 = (b0_4_fu_316_p1 ^ b0_30_fu_1398_p3);

assign b0_18_fu_1632_p2 = (b0_19_fu_1604_p3 ^ b0_17_fu_1526_p2);

assign b0_19_fu_1604_p3 = b0_15_fu_1464_p2[32'd2];

assign b0_1_fu_230_p1 = b[7:0];

assign b0_20_fu_1872_p2 = (b0_24_fu_1840_p4 ^ b0_16_fu_1496_p2);

assign b0_21_fu_1902_p2 = (b0_25_fu_1832_p3 ^ b0_17_fu_1526_p2);

assign b0_22_fu_2008_p2 = (b0_23_fu_1980_p3 ^ b0_21_fu_1902_p2);

assign b0_23_fu_1980_p3 = b_56_fu_1850_p2[32'd2];

assign b0_24_fu_1840_p4 = {{b_42_fu_1436_p2[5:4]}};

assign b0_25_fu_1832_p3 = b_42_fu_1436_p2[32'd4];

assign b0_26_fu_2312_p2 = (b0_27_fu_2284_p3 ^ b0_25_fu_1832_p3);

assign b0_27_fu_2284_p3 = b_42_fu_1436_p2[32'd6];

assign b0_28_fu_1416_p4 = {{b[11:8]}};

assign b0_29_fu_1406_p4 = {{b[9:8]}};

assign b0_2_fu_262_p1 = b[3:0];

assign b0_30_fu_1398_p3 = b[32'd8];

assign b0_31_fu_2708_p2 = (b0_32_fu_2680_p3 ^ b0_30_fu_1398_p3);

assign b0_32_fu_2680_p3 = b[32'd10];

assign b0_33_fu_2948_p2 = (b0_37_fu_2916_p4 ^ b0_29_fu_1406_p4);

assign b0_34_fu_2978_p2 = (b0_38_fu_2908_p3 ^ b0_30_fu_1398_p3);

assign b0_35_fu_3084_p2 = (b0_36_fu_3056_p3 ^ b0_34_fu_2978_p2);

assign b0_36_fu_3056_p3 = b_96_fu_2926_p2[32'd2];

assign b0_37_fu_2916_p4 = {{b[13:12]}};

assign b0_38_fu_2908_p3 = b[32'd12];

assign b0_39_fu_3388_p2 = (b0_40_fu_3360_p3 ^ b0_38_fu_2908_p3);

assign b0_3_fu_290_p1 = b[1:0];

assign b0_40_fu_3360_p3 = b[32'd14];

assign b0_41_fu_3966_p2 = (b0_81_fu_3860_p4 ^ b0_1_fu_230_p1);

assign b0_42_fu_4004_p2 = (b0_82_fu_3850_p4 ^ b0_2_fu_262_p1);

assign b0_43_fu_4036_p2 = (b0_83_fu_3840_p4 ^ b0_3_fu_290_p1);

assign b0_44_fu_4066_p2 = (b0_84_fu_3832_p3 ^ b0_4_fu_316_p1);

assign b0_45_fu_4172_p2 = (b0_46_fu_4144_p3 ^ b0_44_fu_4066_p2);

assign b0_46_fu_4144_p3 = b0_42_fu_4004_p2[32'd2];

assign b0_47_fu_4412_p2 = (b0_51_fu_4380_p4 ^ b0_43_fu_4036_p2);

assign b0_48_fu_4442_p2 = (b0_52_fu_4372_p3 ^ b0_44_fu_4066_p2);

assign b0_49_fu_4548_p2 = (b0_50_fu_4520_p3 ^ b0_48_fu_4442_p2);

assign b0_4_fu_316_p1 = b[0:0];

assign b0_50_fu_4520_p3 = b_137_fu_4390_p2[32'd2];

assign b0_51_fu_4380_p4 = {{b0_41_fu_3966_p2[5:4]}};

assign b0_52_fu_4372_p3 = b0_41_fu_3966_p2[32'd4];

assign b0_53_fu_4852_p2 = (b0_54_fu_4824_p3 ^ b0_52_fu_4372_p3);

assign b0_54_fu_4824_p3 = b0_41_fu_3966_p2[32'd6];

assign b0_55_fu_5216_p2 = (b0_68_fu_5168_p4 ^ b0_42_fu_4004_p2);

assign b0_56_fu_5248_p2 = (b0_69_fu_5158_p4 ^ b0_43_fu_4036_p2);

assign b0_57_fu_5278_p2 = (b0_70_fu_5150_p3 ^ b0_44_fu_4066_p2);

assign b0_58_fu_5384_p2 = (b0_59_fu_5356_p3 ^ b0_57_fu_5278_p2);

assign b0_59_fu_5356_p3 = b0_55_fu_5216_p2[32'd2];

assign b0_5_fu_420_p2 = (b0_6_fu_392_p3 ^ b0_4_fu_316_p1);

assign b0_60_fu_5624_p2 = (b0_64_fu_5592_p4 ^ b0_56_fu_5248_p2);

assign b0_61_fu_5654_p2 = (b0_65_fu_5584_p3 ^ b0_57_fu_5278_p2);

assign b0_62_fu_5760_p2 = (b0_63_fu_5732_p3 ^ b0_61_fu_5654_p2);

assign b0_63_fu_5732_p3 = b_177_fu_5602_p2[32'd2];

assign b0_64_fu_5592_p4 = {{b_163_fu_5188_p2[5:4]}};

assign b0_65_fu_5584_p3 = b_163_fu_5188_p2[32'd4];

assign b0_66_fu_6064_p2 = (b0_67_fu_6036_p3 ^ b0_65_fu_5584_p3);

assign b0_67_fu_6036_p3 = b_163_fu_5188_p2[32'd6];

assign b0_68_fu_5168_p4 = {{b_122_fu_3900_p2[11:8]}};

assign b0_69_fu_5158_p4 = {{b_122_fu_3900_p2[9:8]}};

assign b0_6_fu_392_p3 = b[32'd2];

assign b0_70_fu_5150_p3 = b_122_fu_3900_p2[32'd8];

assign b0_71_fu_6460_p2 = (b0_72_fu_6432_p3 ^ b0_70_fu_5150_p3);

assign b0_72_fu_6432_p3 = xor_ln33_3_fu_3918_p2[32'd10];

assign b0_73_fu_6700_p2 = (b0_77_fu_6668_p4 ^ b0_69_fu_5158_p4);

assign b0_74_fu_6730_p2 = (b0_78_fu_6660_p3 ^ b0_70_fu_5150_p3);

assign b0_75_fu_6836_p2 = (b0_76_fu_6808_p3 ^ b0_74_fu_6730_p2);

assign b0_76_fu_6808_p3 = b_217_fu_6678_p2[32'd2];

assign b0_77_fu_6668_p4 = {{b_122_fu_3900_p2[13:12]}};

assign b0_78_fu_6660_p3 = b_122_fu_3900_p2[32'd12];

assign b0_79_fu_7140_p2 = (b0_80_fu_7112_p3 ^ b0_78_fu_6660_p3);

assign b0_7_fu_660_p2 = (b0_3_fu_290_p1 ^ b0_11_fu_628_p4);

assign b0_80_fu_7112_p3 = b_122_fu_3900_p2[32'd14];

assign b0_81_fu_3860_p4 = {{b[23:16]}};

assign b0_82_fu_3850_p4 = {{b[19:16]}};

assign b0_83_fu_3840_p4 = {{b[17:16]}};

assign b0_84_fu_3832_p3 = b[32'd16];

assign b0_85_fu_7660_p2 = (b0_86_fu_7632_p3 ^ b0_84_fu_3832_p3);

assign b0_86_fu_7632_p3 = b[32'd18];

assign b0_87_fu_7900_p2 = (b0_91_fu_7868_p4 ^ b0_83_fu_3840_p4);

assign b0_88_fu_7930_p2 = (b0_92_fu_7860_p3 ^ b0_84_fu_3832_p3);

assign b0_89_fu_8036_p2 = (b0_90_fu_8008_p3 ^ b0_88_fu_7930_p2);

assign b0_8_fu_690_p2 = (b0_4_fu_316_p1 ^ b0_12_fu_620_p3);

assign b0_90_fu_8008_p3 = b_258_fu_7878_p2[32'd2];

assign b0_91_fu_7868_p4 = {{b[21:20]}};

assign b0_92_fu_7860_p3 = b[32'd20];

assign b0_93_fu_8340_p2 = (b0_94_fu_8312_p3 ^ b0_92_fu_7860_p3);

assign b0_94_fu_8312_p3 = b[32'd22];

assign b0_95_fu_8704_p2 = (b0_82_fu_3850_p4 ^ b0_108_fu_8656_p4);

assign b0_96_fu_8736_p2 = (b0_83_fu_3840_p4 ^ b0_109_fu_8646_p4);

assign b0_97_fu_8766_p2 = (b0_84_fu_3832_p3 ^ b0_110_fu_8638_p3);

assign b0_98_fu_8872_p2 = (b0_99_fu_8844_p3 ^ b0_97_fu_8766_p2);

assign b0_99_fu_8844_p3 = b0_95_fu_8704_p2[32'd2];

assign b0_9_fu_796_p2 = (b0_8_fu_690_p2 ^ b0_10_fu_768_p3);

assign b0_fu_186_p1 = b[15:0];

assign b1_117_fu_238_p4 = {{b[15:8]}};

assign b1_118_fu_266_p4 = {{b[7:4]}};

assign b1_119_fu_294_p4 = {{b[3:2]}};

assign b1_120_fu_320_p3 = b[32'd1];

assign b1_121_fu_426_p3 = b_8_fu_400_p2[32'd1];

assign b1_122_fu_492_p3 = b[32'd3];

assign b1_123_fu_666_p4 = {{b_16_fu_638_p2[3:2]}};

assign b1_124_fu_696_p3 = b0_7_fu_660_p2[32'd1];

assign b1_125_fu_802_p3 = b_21_fu_776_p2[32'd1];

assign b1_126_fu_868_p3 = b_16_fu_638_p2[32'd3];

assign b1_127_fu_982_p4 = {{b[7:6]}};

assign b1_128_fu_1000_p3 = b[32'd5];

assign b1_129_fu_1106_p3 = b_34_fu_1080_p2[32'd1];

assign b1_130_fu_1172_p3 = b[32'd7];

assign b1_131_fu_1470_p4 = {{b_42_fu_1436_p2[7:4]}};

assign b1_132_fu_1502_p4 = {{b0_15_fu_1464_p2[3:2]}};

assign b1_133_fu_1532_p3 = b0_16_fu_1496_p2[32'd1];

assign b1_134_fu_1638_p3 = b_48_fu_1612_p2[32'd1];

assign b1_135_fu_1704_p3 = b0_15_fu_1464_p2[32'd3];

assign b1_136_fu_1878_p4 = {{b_56_fu_1850_p2[3:2]}};

assign b1_137_fu_1908_p3 = b0_20_fu_1872_p2[32'd1];

assign b1_138_fu_2014_p3 = b_61_fu_1988_p2[32'd1];

assign b1_139_fu_2080_p3 = b_56_fu_1850_p2[32'd3];

assign b1_140_fu_2194_p4 = {{b_42_fu_1436_p2[7:6]}};

assign b1_141_fu_2212_p3 = xor_ln33_fu_1442_p2[32'd5];

assign b1_142_fu_2318_p3 = b_74_fu_2292_p2[32'd1];

assign b1_143_fu_2384_p3 = b_42_fu_1436_p2[32'd7];

assign b1_144_fu_2570_p4 = {{b[15:12]}};

assign b1_145_fu_2590_p4 = {{b[11:10]}};

assign b1_146_fu_2608_p3 = b[32'd9];

assign b1_147_fu_2714_p3 = b_88_fu_2688_p2[32'd1];

assign b1_148_fu_2780_p3 = b[32'd11];

assign b1_149_fu_2954_p4 = {{b_96_fu_2926_p2[3:2]}};

assign b1_150_fu_2984_p3 = b0_33_fu_2948_p2[32'd1];

assign b1_151_fu_3090_p3 = b_101_fu_3064_p2[32'd1];

assign b1_152_fu_3156_p3 = b_96_fu_2926_p2[32'd3];

assign b1_153_fu_3270_p4 = {{b[15:14]}};

assign b1_154_fu_3288_p3 = b[32'd13];

assign b1_155_fu_3394_p3 = b_114_fu_3368_p2[32'd1];

assign b1_156_fu_3460_p3 = b[32'd15];

assign b1_157_fu_3978_p4 = {{b_122_fu_3900_p2[15:8]}};

assign b1_158_fu_4010_p4 = {{b0_41_fu_3966_p2[7:4]}};

assign b1_159_fu_4042_p4 = {{b0_42_fu_4004_p2[3:2]}};

assign b1_160_fu_4072_p3 = b0_43_fu_4036_p2[32'd1];

assign b1_161_fu_4178_p3 = b_129_fu_4152_p2[32'd1];

assign b1_162_fu_4244_p3 = b0_42_fu_4004_p2[32'd3];

assign b1_163_fu_4418_p4 = {{b_137_fu_4390_p2[3:2]}};

assign b1_164_fu_4448_p3 = b0_47_fu_4412_p2[32'd1];

assign b1_165_fu_4554_p3 = b_142_fu_4528_p2[32'd1];

assign b1_166_fu_4620_p3 = b_137_fu_4390_p2[32'd3];

assign b1_167_fu_4734_p4 = {{b0_41_fu_3966_p2[7:6]}};

assign b1_168_fu_4752_p3 = xor_ln40_1_fu_3972_p2[32'd5];

assign b1_169_fu_4858_p3 = b_155_fu_4832_p2[32'd1];

assign b1_170_fu_4924_p3 = b0_41_fu_3966_p2[32'd7];

assign b1_171_fu_5222_p4 = {{b_163_fu_5188_p2[7:4]}};

assign b1_172_fu_5254_p4 = {{b0_55_fu_5216_p2[3:2]}};

assign b1_173_fu_5284_p3 = b0_56_fu_5248_p2[32'd1];

assign b1_174_fu_5390_p3 = b_169_fu_5364_p2[32'd1];

assign b1_175_fu_5456_p3 = b0_55_fu_5216_p2[32'd3];

assign b1_176_fu_5630_p4 = {{b_177_fu_5602_p2[3:2]}};

assign b1_177_fu_5660_p3 = b0_60_fu_5624_p2[32'd1];

assign b1_178_fu_5766_p3 = b_182_fu_5740_p2[32'd1];

assign b1_179_fu_5832_p3 = b_177_fu_5602_p2[32'd3];

assign b1_180_fu_5946_p4 = {{b_163_fu_5188_p2[7:6]}};

assign b1_181_fu_5964_p3 = xor_ln33_4_fu_5194_p2[32'd5];

assign b1_182_fu_6070_p3 = b_195_fu_6044_p2[32'd1];

assign b1_183_fu_6136_p3 = b_163_fu_5188_p2[32'd7];

assign b1_184_fu_6322_p4 = {{b_122_fu_3900_p2[15:12]}};

assign b1_185_fu_6342_p4 = {{xor_ln33_3_fu_3918_p2[11:10]}};

assign b1_186_fu_6360_p3 = xor_ln33_2_fu_3912_p2[32'd9];

assign b1_187_fu_6466_p3 = b_209_fu_6440_p2[32'd1];

assign b1_188_fu_6532_p3 = xor_ln33_3_fu_3918_p2[32'd11];

assign b1_189_fu_6706_p4 = {{b_217_fu_6678_p2[3:2]}};

assign b1_190_fu_6736_p3 = b0_73_fu_6700_p2[32'd1];

assign b1_191_fu_6842_p3 = b_222_fu_6816_p2[32'd1];

assign b1_192_fu_6908_p3 = b_217_fu_6678_p2[32'd3];

assign b1_193_fu_7022_p4 = {{b_122_fu_3900_p2[15:14]}};

assign b1_194_fu_7040_p3 = xor_ln33_1_fu_3906_p2[32'd13];

assign b1_195_fu_7146_p3 = b_235_fu_7120_p2[32'd1];

assign b1_196_fu_7212_p3 = b_122_fu_3900_p2[32'd15];

assign b1_197_fu_7502_p4 = {{b[31:24]}};

assign b1_198_fu_7522_p4 = {{b[23:20]}};

assign b1_199_fu_7542_p4 = {{b[19:18]}};

assign b1_200_fu_7560_p3 = b[32'd17];

assign b1_201_fu_7666_p3 = b_250_fu_7640_p2[32'd1];

assign b1_202_fu_7732_p3 = b[32'd19];

assign b1_203_fu_7906_p4 = {{b_258_fu_7878_p2[3:2]}};

assign b1_204_fu_7936_p3 = b0_87_fu_7900_p2[32'd1];

assign b1_205_fu_8042_p3 = b_263_fu_8016_p2[32'd1];

assign b1_206_fu_8108_p3 = b_258_fu_7878_p2[32'd3];

assign b1_207_fu_8222_p4 = {{b[23:22]}};

assign b1_208_fu_8240_p3 = b[32'd21];

assign b1_209_fu_8346_p3 = b_276_fu_8320_p2[32'd1];

assign b1_210_fu_8412_p3 = b[32'd23];

assign b1_211_fu_8710_p4 = {{b_284_fu_8676_p2[7:4]}};

assign b1_212_fu_8742_p4 = {{b0_95_fu_8704_p2[3:2]}};

assign b1_213_fu_8772_p3 = b0_96_fu_8736_p2[32'd1];

assign b1_214_fu_8878_p3 = b_290_fu_8852_p2[32'd1];

assign b1_215_fu_8944_p3 = b0_95_fu_8704_p2[32'd3];

assign b1_216_fu_9118_p4 = {{b_298_fu_9090_p2[3:2]}};

assign b1_217_fu_9148_p3 = b0_100_fu_9112_p2[32'd1];

assign b1_218_fu_9254_p3 = b_303_fu_9228_p2[32'd1];

assign b1_219_fu_9320_p3 = b_298_fu_9090_p2[32'd3];

assign b1_220_fu_9434_p4 = {{b_284_fu_8676_p2[7:6]}};

assign b1_221_fu_9452_p3 = xor_ln33_5_fu_8682_p2[32'd5];

assign b1_222_fu_9558_p3 = b_316_fu_9532_p2[32'd1];

assign b1_223_fu_9624_p3 = b_284_fu_8676_p2[32'd7];

assign b1_224_fu_9810_p4 = {{b[31:28]}};

assign b1_225_fu_9830_p4 = {{b[27:26]}};

assign b1_226_fu_9848_p3 = b[32'd25];

assign b1_227_fu_9954_p3 = b_330_fu_9928_p2[32'd1];

assign b1_228_fu_10020_p3 = b[32'd27];

assign b1_229_fu_10194_p4 = {{b_338_fu_10166_p2[3:2]}};

assign b1_230_fu_10224_p3 = b0_113_fu_10188_p2[32'd1];

assign b1_231_fu_10330_p3 = b_343_fu_10304_p2[32'd1];

assign b1_232_fu_10396_p3 = b_338_fu_10166_p2[32'd3];

assign b1_233_fu_10510_p4 = {{b[31:30]}};

assign b1_234_fu_10528_p3 = b[32'd29];

assign b1_235_fu_10634_p3 = b_356_fu_10608_p2[32'd1];

assign b1_236_fu_10700_p3 = b[32'd31];

assign b1_fu_202_p4 = {{b[31:16]}};

assign b_101_fu_3064_p2 = (b1_149_fu_2954_p4 ^ b0_33_fu_2948_p2);

assign b_103_fu_3110_p2 = (b1_151_fu_3090_p3 ^ b0_35_fu_3084_p2);

assign b_107_fu_3176_p2 = (b1_152_fu_3156_p3 ^ b0_36_fu_3056_p3);

assign b_10_fu_446_p2 = (b1_121_fu_426_p3 ^ b0_5_fu_420_p2);

assign b_112_fu_3308_p2 = (b1_154_fu_3288_p3 ^ b0_38_fu_2908_p3);

assign b_114_fu_3368_p2 = (b1_153_fu_3270_p4 ^ b0_37_fu_2916_p4);

assign b_116_fu_3414_p2 = (b1_155_fu_3394_p3 ^ b0_39_fu_3388_p2);

assign b_120_fu_3480_p2 = (b1_156_fu_3460_p3 ^ b0_40_fu_3360_p3);

assign b_122_fu_3900_p2 = (b1_fu_202_p4 ^ b0_fu_186_p1);

assign b_127_fu_4092_p2 = (b1_160_fu_4072_p3 ^ b0_44_fu_4066_p2);

assign b_129_fu_4152_p2 = (b1_159_fu_4042_p4 ^ b0_43_fu_4036_p2);

assign b_131_fu_4198_p2 = (b1_161_fu_4178_p3 ^ b0_45_fu_4172_p2);

assign b_135_fu_4264_p2 = (b1_162_fu_4244_p3 ^ b0_46_fu_4144_p3);

assign b_137_fu_4390_p2 = (b1_158_fu_4010_p4 ^ b0_42_fu_4004_p2);

assign b_140_fu_4468_p2 = (b1_164_fu_4448_p3 ^ b0_48_fu_4442_p2);

assign b_142_fu_4528_p2 = (b1_163_fu_4418_p4 ^ b0_47_fu_4412_p2);

assign b_144_fu_4574_p2 = (b1_165_fu_4554_p3 ^ b0_49_fu_4548_p2);

assign b_148_fu_4640_p2 = (b1_166_fu_4620_p3 ^ b0_50_fu_4520_p3);

assign b_14_fu_512_p2 = (b1_122_fu_492_p3 ^ b0_6_fu_392_p3);

assign b_153_fu_4772_p2 = (b1_168_fu_4752_p3 ^ b0_52_fu_4372_p3);

assign b_155_fu_4832_p2 = (b1_167_fu_4734_p4 ^ b0_51_fu_4380_p4);

assign b_157_fu_4878_p2 = (b1_169_fu_4858_p3 ^ b0_53_fu_4852_p2);

assign b_161_fu_4944_p2 = (b1_170_fu_4924_p3 ^ b0_54_fu_4824_p3);

assign b_163_fu_5188_p2 = (b1_157_fu_3978_p4 ^ b0_41_fu_3966_p2);

assign b_167_fu_5304_p2 = (b1_173_fu_5284_p3 ^ b0_57_fu_5278_p2);

assign b_169_fu_5364_p2 = (b1_172_fu_5254_p4 ^ b0_56_fu_5248_p2);

assign b_16_fu_638_p2 = (b1_118_fu_266_p4 ^ b0_2_fu_262_p1);

assign b_171_fu_5410_p2 = (b1_174_fu_5390_p3 ^ b0_58_fu_5384_p2);

assign b_175_fu_5476_p2 = (b1_175_fu_5456_p3 ^ b0_59_fu_5356_p3);

assign b_177_fu_5602_p2 = (b1_171_fu_5222_p4 ^ b0_55_fu_5216_p2);

assign b_180_fu_5680_p2 = (b1_177_fu_5660_p3 ^ b0_61_fu_5654_p2);

assign b_182_fu_5740_p2 = (b1_176_fu_5630_p4 ^ b0_60_fu_5624_p2);

assign b_184_fu_5786_p2 = (b1_178_fu_5766_p3 ^ b0_62_fu_5760_p2);

assign b_188_fu_5852_p2 = (b1_179_fu_5832_p3 ^ b0_63_fu_5732_p3);

assign b_193_fu_5984_p2 = (b1_181_fu_5964_p3 ^ b0_65_fu_5584_p3);

assign b_195_fu_6044_p2 = (b1_180_fu_5946_p4 ^ b0_64_fu_5592_p4);

assign b_197_fu_6090_p2 = (b1_182_fu_6070_p3 ^ b0_66_fu_6064_p2);

assign b_19_fu_716_p2 = (b1_124_fu_696_p3 ^ b0_8_fu_690_p2);

assign b_201_fu_6156_p2 = (b1_183_fu_6136_p3 ^ b0_67_fu_6036_p3);

assign b_207_fu_6380_p2 = (b1_186_fu_6360_p3 ^ b0_70_fu_5150_p3);

assign b_209_fu_6440_p2 = (b1_185_fu_6342_p4 ^ b0_69_fu_5158_p4);

assign b_211_fu_6486_p2 = (b1_187_fu_6466_p3 ^ b0_71_fu_6460_p2);

assign b_215_fu_6552_p2 = (b1_188_fu_6532_p3 ^ b0_72_fu_6432_p3);

assign b_217_fu_6678_p2 = (b1_184_fu_6322_p4 ^ b0_68_fu_5168_p4);

assign b_21_fu_776_p2 = (b1_123_fu_666_p4 ^ b0_7_fu_660_p2);

assign b_220_fu_6756_p2 = (b1_190_fu_6736_p3 ^ b0_74_fu_6730_p2);

assign b_222_fu_6816_p2 = (b1_189_fu_6706_p4 ^ b0_73_fu_6700_p2);

assign b_224_fu_6862_p2 = (b1_191_fu_6842_p3 ^ b0_75_fu_6836_p2);

assign b_228_fu_6928_p2 = (b1_192_fu_6908_p3 ^ b0_76_fu_6808_p3);

assign b_233_fu_7060_p2 = (b1_194_fu_7040_p3 ^ b0_78_fu_6660_p3);

assign b_235_fu_7120_p2 = (b1_193_fu_7022_p4 ^ b0_77_fu_6668_p4);

assign b_237_fu_7166_p2 = (b1_195_fu_7146_p3 ^ b0_79_fu_7140_p2);

assign b_23_fu_822_p2 = (b1_125_fu_802_p3 ^ b0_9_fu_796_p2);

assign b_241_fu_7232_p2 = (b1_196_fu_7212_p3 ^ b0_80_fu_7112_p3);

assign b_248_fu_7580_p2 = (b1_200_fu_7560_p3 ^ b0_84_fu_3832_p3);

assign b_250_fu_7640_p2 = (b1_199_fu_7542_p4 ^ b0_83_fu_3840_p4);

assign b_252_fu_7686_p2 = (b1_201_fu_7666_p3 ^ b0_85_fu_7660_p2);

assign b_256_fu_7752_p2 = (b1_202_fu_7732_p3 ^ b0_86_fu_7632_p3);

assign b_258_fu_7878_p2 = (b1_198_fu_7522_p4 ^ b0_82_fu_3850_p4);

assign b_261_fu_7956_p2 = (b1_204_fu_7936_p3 ^ b0_88_fu_7930_p2);

assign b_263_fu_8016_p2 = (b1_203_fu_7906_p4 ^ b0_87_fu_7900_p2);

assign b_265_fu_8062_p2 = (b1_205_fu_8042_p3 ^ b0_89_fu_8036_p2);

assign b_269_fu_8128_p2 = (b1_206_fu_8108_p3 ^ b0_90_fu_8008_p3);

assign b_274_fu_8260_p2 = (b1_208_fu_8240_p3 ^ b0_92_fu_7860_p3);

assign b_276_fu_8320_p2 = (b1_207_fu_8222_p4 ^ b0_91_fu_7868_p4);

assign b_278_fu_8366_p2 = (b1_209_fu_8346_p3 ^ b0_93_fu_8340_p2);

assign b_27_fu_888_p2 = (b1_126_fu_868_p3 ^ b0_10_fu_768_p3);

assign b_282_fu_8432_p2 = (b1_210_fu_8412_p3 ^ b0_94_fu_8312_p3);

assign b_284_fu_8676_p2 = (b1_197_fu_7502_p4 ^ b0_81_fu_3860_p4);

assign b_288_fu_8792_p2 = (b1_213_fu_8772_p3 ^ b0_97_fu_8766_p2);

assign b_290_fu_8852_p2 = (b1_212_fu_8742_p4 ^ b0_96_fu_8736_p2);

assign b_292_fu_8898_p2 = (b1_214_fu_8878_p3 ^ b0_98_fu_8872_p2);

assign b_296_fu_8964_p2 = (b1_215_fu_8944_p3 ^ b0_99_fu_8844_p3);

assign b_298_fu_9090_p2 = (b1_211_fu_8710_p4 ^ b0_95_fu_8704_p2);

assign b_301_fu_9168_p2 = (b1_217_fu_9148_p3 ^ b0_101_fu_9142_p2);

assign b_303_fu_9228_p2 = (b1_216_fu_9118_p4 ^ b0_100_fu_9112_p2);

assign b_305_fu_9274_p2 = (b1_218_fu_9254_p3 ^ b0_102_fu_9248_p2);

assign b_309_fu_9340_p2 = (b1_219_fu_9320_p3 ^ b0_103_fu_9220_p3);

assign b_314_fu_9472_p2 = (b1_221_fu_9452_p3 ^ b0_105_fu_9072_p3);

assign b_316_fu_9532_p2 = (b1_220_fu_9434_p4 ^ b0_104_fu_9080_p4);

assign b_318_fu_9578_p2 = (b1_222_fu_9558_p3 ^ b0_106_fu_9552_p2);

assign b_322_fu_9644_p2 = (b1_223_fu_9624_p3 ^ b0_107_fu_9524_p3);

assign b_328_fu_9868_p2 = (b1_226_fu_9848_p3 ^ b0_110_fu_8638_p3);

assign b_32_fu_1020_p2 = (b1_128_fu_1000_p3 ^ b0_12_fu_620_p3);

assign b_330_fu_9928_p2 = (b1_225_fu_9830_p4 ^ b0_109_fu_8646_p4);

assign b_332_fu_9974_p2 = (b1_227_fu_9954_p3 ^ b0_111_fu_9948_p2);

assign b_336_fu_10040_p2 = (b1_228_fu_10020_p3 ^ b0_112_fu_9920_p3);

assign b_338_fu_10166_p2 = (b1_224_fu_9810_p4 ^ b0_108_fu_8656_p4);

assign b_341_fu_10244_p2 = (b1_230_fu_10224_p3 ^ b0_114_fu_10218_p2);

assign b_343_fu_10304_p2 = (b1_229_fu_10194_p4 ^ b0_113_fu_10188_p2);

assign b_345_fu_10350_p2 = (b1_231_fu_10330_p3 ^ b0_115_fu_10324_p2);

assign b_349_fu_10416_p2 = (b1_232_fu_10396_p3 ^ b0_116_fu_10296_p3);

assign b_34_fu_1080_p2 = (b1_127_fu_982_p4 ^ b0_11_fu_628_p4);

assign b_354_fu_10548_p2 = (b1_234_fu_10528_p3 ^ b0_118_fu_10148_p3);

assign b_356_fu_10608_p2 = (b1_233_fu_10510_p4 ^ b0_117_fu_10156_p4);

assign b_358_fu_10654_p2 = (b1_235_fu_10634_p3 ^ b0_119_fu_10628_p2);

assign b_362_fu_10720_p2 = (b1_236_fu_10700_p3 ^ b0_120_fu_10600_p3);

assign b_36_fu_1126_p2 = (b1_129_fu_1106_p3 ^ b0_13_fu_1100_p2);

assign b_40_fu_1192_p2 = (b1_130_fu_1172_p3 ^ b0_14_fu_1072_p3);

assign b_42_fu_1436_p2 = (b1_117_fu_238_p4 ^ b0_1_fu_230_p1);

assign b_46_fu_1552_p2 = (b1_133_fu_1532_p3 ^ b0_17_fu_1526_p2);

assign b_48_fu_1612_p2 = (b1_132_fu_1502_p4 ^ b0_16_fu_1496_p2);

assign b_50_fu_1658_p2 = (b1_134_fu_1638_p3 ^ b0_18_fu_1632_p2);

assign b_54_fu_1724_p2 = (b1_135_fu_1704_p3 ^ b0_19_fu_1604_p3);

assign b_56_fu_1850_p2 = (b1_131_fu_1470_p4 ^ b0_15_fu_1464_p2);

assign b_59_fu_1928_p2 = (b1_137_fu_1908_p3 ^ b0_21_fu_1902_p2);

assign b_61_fu_1988_p2 = (b1_136_fu_1878_p4 ^ b0_20_fu_1872_p2);

assign b_63_fu_2034_p2 = (b1_138_fu_2014_p3 ^ b0_22_fu_2008_p2);

assign b_67_fu_2100_p2 = (b1_139_fu_2080_p3 ^ b0_23_fu_1980_p3);

assign b_6_fu_340_p2 = (b1_120_fu_320_p3 ^ b0_4_fu_316_p1);

assign b_72_fu_2232_p2 = (b1_141_fu_2212_p3 ^ b0_25_fu_1832_p3);

assign b_74_fu_2292_p2 = (b1_140_fu_2194_p4 ^ b0_24_fu_1840_p4);

assign b_76_fu_2338_p2 = (b1_142_fu_2318_p3 ^ b0_26_fu_2312_p2);

assign b_80_fu_2404_p2 = (b1_143_fu_2384_p3 ^ b0_27_fu_2284_p3);

assign b_86_fu_2628_p2 = (b1_146_fu_2608_p3 ^ b0_30_fu_1398_p3);

assign b_88_fu_2688_p2 = (b1_145_fu_2590_p4 ^ b0_29_fu_1406_p4);

assign b_8_fu_400_p2 = (b1_119_fu_294_p4 ^ b0_3_fu_290_p1);

assign b_90_fu_2734_p2 = (b1_147_fu_2714_p3 ^ b0_31_fu_2708_p2);

assign b_94_fu_2800_p2 = (b1_148_fu_2780_p3 ^ b0_32_fu_2680_p3);

assign b_96_fu_2926_p2 = (b1_144_fu_2570_p4 ^ b0_28_fu_1416_p4);

assign b_99_fu_3004_p2 = (b1_150_fu_2984_p3 ^ b0_34_fu_2978_p2);

assign tmp_10_fu_3220_p3 = {{xor_ln28_11_fu_3214_p2}, {a1_58_fu_3194_p2}};

assign tmp_11_fu_3524_p3 = {{xor_ln28_12_fu_3518_p2}, {a1_63_fu_3498_p2}};

assign tmp_12_fu_3582_p3 = {{xor_ln28_13_fu_3576_p2}, {a1_66_fu_3568_p3}};

assign tmp_13_fu_3596_p3 = {{xor_ln28_14_fu_3590_p2}, {a1_248_fu_3544_p2}};

assign tmp_14_fu_3672_p3 = {{xor_ln28_15_fu_3666_p2}, {a1_69_fu_3658_p3}};

assign tmp_15_fu_3686_p3 = {{xor_ln28_16_fu_3680_p2}, {a1_250_fu_3640_p4}};

assign tmp_16_fu_3700_p3 = {{xor_ln28_17_fu_3694_p2}, {a1_249_fu_3616_p2}};

assign tmp_17_fu_4308_p3 = {{xor_ln28_18_fu_4302_p2}, {a1_78_fu_4282_p2}};

assign tmp_18_fu_4684_p3 = {{xor_ln28_19_fu_4678_p2}, {a1_84_fu_4658_p2}};

assign tmp_19_fu_4988_p3 = {{xor_ln28_20_fu_4982_p2}, {a1_90_fu_4962_p2}};

assign tmp_1_fu_1294_p3 = {{xor_ln28_3_fu_1288_p2}, {a1_23_fu_1280_p3}};

assign tmp_20_fu_5046_p3 = {{xor_ln28_21_fu_5040_p2}, {a1_92_fu_5032_p3}};

assign tmp_21_fu_5060_p3 = {{xor_ln28_22_fu_5054_p2}, {a1_265_fu_5008_p2}};

assign tmp_22_fu_5520_p3 = {{xor_ln28_23_fu_5514_p2}, {a1_99_fu_5494_p2}};

assign tmp_23_fu_5896_p3 = {{xor_ln28_24_fu_5890_p2}, {a1_105_fu_5870_p2}};

assign tmp_24_fu_6200_p3 = {{xor_ln28_25_fu_6194_p2}, {a1_112_fu_6174_p2}};

assign tmp_25_fu_6258_p3 = {{xor_ln28_26_fu_6252_p2}, {a1_114_fu_6244_p3}};

assign tmp_26_fu_6272_p3 = {{xor_ln28_27_fu_6266_p2}, {a1_279_fu_6220_p2}};

assign tmp_27_fu_6596_p3 = {{xor_ln28_28_fu_6590_p2}, {a1_120_fu_6570_p2}};

assign tmp_28_fu_6972_p3 = {{xor_ln28_29_fu_6966_p2}, {a1_126_fu_6946_p2}};

assign tmp_29_fu_7276_p3 = {{xor_ln28_30_fu_7270_p2}, {a1_133_fu_7250_p2}};

assign tmp_2_fu_1308_p3 = {{xor_ln28_4_fu_1302_p2}, {a1_220_fu_1256_p2}};

assign tmp_30_fu_7334_p3 = {{xor_ln28_31_fu_7328_p2}, {a1_135_fu_7320_p3}};

assign tmp_31_fu_7348_p3 = {{xor_ln28_32_fu_7342_p2}, {a1_293_fu_7296_p2}};

assign tmp_32_fu_7424_p3 = {{xor_ln28_33_fu_7418_p2}, {a1_138_fu_7410_p3}};

assign tmp_33_fu_7438_p3 = {{xor_ln28_34_fu_7432_p2}, {a1_295_fu_7392_p4}};

assign tmp_34_fu_7452_p3 = {{xor_ln28_35_fu_7446_p2}, {a1_294_fu_7368_p2}};

assign tmp_35_fu_7796_p3 = {{xor_ln28_36_fu_7790_p2}, {a1_147_fu_7770_p2}};

assign tmp_36_fu_8172_p3 = {{xor_ln28_37_fu_8166_p2}, {a1_153_fu_8146_p2}};

assign tmp_37_fu_8476_p3 = {{xor_ln28_38_fu_8470_p2}, {a1_159_fu_8450_p2}};

assign tmp_38_fu_8534_p3 = {{xor_ln28_39_fu_8528_p2}, {a1_161_fu_8520_p3}};

assign tmp_39_fu_8548_p3 = {{xor_ln28_40_fu_8542_p2}, {a1_310_fu_8496_p2}};

assign tmp_3_fu_1768_p3 = {{xor_ln28_5_fu_1762_p2}, {a1_31_fu_1742_p2}};

assign tmp_40_fu_9008_p3 = {{xor_ln28_41_fu_9002_p2}, {a1_168_fu_8982_p2}};

assign tmp_41_fu_9384_p3 = {{xor_ln28_42_fu_9378_p2}, {a1_173_fu_9358_p2}};

assign tmp_42_fu_9688_p3 = {{xor_ln28_43_fu_9682_p2}, {a1_178_fu_9662_p2}};

assign tmp_43_fu_9746_p3 = {{xor_ln28_44_fu_9740_p2}, {a1_180_fu_9732_p3}};

assign tmp_44_fu_9760_p3 = {{xor_ln28_45_fu_9754_p2}, {a1_324_fu_9708_p2}};

assign tmp_45_fu_10084_p3 = {{xor_ln28_46_fu_10078_p2}, {a1_186_fu_10058_p2}};

assign tmp_46_fu_10460_p3 = {{xor_ln28_47_fu_10454_p2}, {a1_191_fu_10434_p2}};

assign tmp_47_fu_10764_p3 = {{xor_ln28_48_fu_10758_p2}, {a1_fu_10738_p2}};

assign tmp_48_fu_10822_p3 = {{xor_ln28_49_fu_10816_p2}, {a1_197_fu_10808_p3}};

assign tmp_49_fu_10836_p3 = {{xor_ln28_50_fu_10830_p2}, {a1_338_fu_10784_p2}};

assign tmp_4_fu_2144_p3 = {{xor_ln28_6_fu_2138_p2}, {a1_37_fu_2118_p2}};

assign tmp_50_fu_10912_p3 = {{xor_ln28_51_fu_10906_p2}, {a1_200_fu_10898_p3}};

assign tmp_51_fu_10926_p3 = {{xor_ln28_52_fu_10920_p2}, {a1_340_fu_10880_p4}};

assign tmp_52_fu_10940_p3 = {{xor_ln28_53_fu_10934_p2}, {a1_339_fu_10856_p2}};

assign tmp_53_fu_11036_p3 = {{xor_ln28_54_fu_11030_p2}, {a1_204_fu_11022_p3}};

assign tmp_54_fu_11050_p3 = {{xor_ln28_55_fu_11044_p2}, {a1_343_fu_11004_p4}};

assign tmp_55_fu_11064_p3 = {{xor_ln28_56_fu_11058_p2}, {a1_342_fu_10984_p4}};

assign tmp_56_fu_11078_p3 = {{xor_ln28_57_fu_11072_p2}, {a1_341_fu_10960_p2}};

assign tmp_5_fu_932_p3 = {{xor_ln28_1_fu_926_p2}, {a1_15_fu_906_p2}};

assign tmp_6_fu_2448_p3 = {{xor_ln28_7_fu_2442_p2}, {a1_42_fu_2422_p2}};

assign tmp_7_fu_2506_p3 = {{xor_ln28_8_fu_2500_p2}, {a1_45_fu_2492_p3}};

assign tmp_8_fu_2520_p3 = {{xor_ln28_9_fu_2514_p2}, {a1_234_fu_2468_p2}};

assign tmp_9_fu_2844_p3 = {{xor_ln28_10_fu_2838_p2}, {a1_52_fu_2818_p2}};

assign tmp_fu_556_p3 = {{xor_ln28_fu_550_p2}, {a1_9_fu_530_p2}};

assign tmp_s_fu_1236_p3 = {{xor_ln28_2_fu_1230_p2}, {a1_21_fu_1210_p2}};

assign trunc_ln38_1_fu_164_p1 = a[13:0];

assign trunc_ln38_2_fu_168_p1 = a[9:0];

assign trunc_ln38_3_fu_172_p1 = a[11:0];

assign trunc_ln38_4_fu_216_p1 = a[5:0];

assign trunc_ln38_5_fu_3924_p4 = {{a[21:16]}};

assign trunc_ln40_1_fu_190_p1 = b[13:0];

assign trunc_ln40_2_fu_194_p1 = b[9:0];

assign trunc_ln40_3_fu_198_p1 = b[11:0];

assign trunc_ln40_4_fu_234_p1 = b[5:0];

assign trunc_ln40_5_fu_3956_p4 = {{b[21:16]}};

assign trunc_ln43_10_fu_8616_p4 = {{a[29:24]}};

assign trunc_ln43_11_fu_8666_p4 = {{b[29:24]}};

assign trunc_ln43_1_fu_1426_p4 = {{b[13:8]}};

assign trunc_ln43_2_fu_3778_p4 = {{a[27:16]}};

assign trunc_ln43_3_fu_3788_p4 = {{a[25:16]}};

assign trunc_ln43_4_fu_3798_p4 = {{a[29:16]}};

assign trunc_ln43_5_fu_3870_p4 = {{b[27:16]}};

assign trunc_ln43_6_fu_3880_p4 = {{b[25:16]}};

assign trunc_ln43_7_fu_3890_p4 = {{b[29:16]}};

assign trunc_ln43_8_fu_5128_p4 = {{a_140_fu_3808_p2[13:8]}};

assign trunc_ln43_9_fu_5178_p4 = {{b_122_fu_3900_p2[13:8]}};

assign trunc_ln43_s_fu_1376_p4 = {{a[13:8]}};

assign xor_ln28_10_fu_2838_p2 = (z2_28_fu_2812_p2 ^ z1_30_fu_2806_p2);

assign xor_ln28_11_fu_3214_p2 = (z2_32_fu_3188_p2 ^ z1_34_fu_3182_p2);

assign xor_ln28_12_fu_3518_p2 = (z2_36_fu_3492_p2 ^ z1_39_fu_3486_p2);

assign xor_ln28_13_fu_3576_p2 = (a1_66_fu_3568_p3 ^ a0_74_fu_3564_p1);

assign xor_ln28_14_fu_3590_p2 = (tmp_12_fu_3582_p3 ^ a0_72_fu_3550_p2);

assign xor_ln28_15_fu_3666_p2 = (a1_69_fu_3658_p3 ^ a0_78_fu_3650_p3);

assign xor_ln28_16_fu_3680_p2 = (tmp_14_fu_3672_p3 ^ a0_76_fu_3636_p1);

assign xor_ln28_17_fu_3694_p2 = (tmp_15_fu_3686_p3 ^ a0_75_fu_3622_p2);

assign xor_ln28_18_fu_4302_p2 = (z2_42_fu_4276_p2 ^ z1_43_fu_4270_p2);

assign xor_ln28_19_fu_4678_p2 = (z2_46_fu_4652_p2 ^ z1_47_fu_4646_p2);

assign xor_ln28_1_fu_926_p2 = (z2_6_fu_900_p2 ^ z1_7_fu_894_p2);

assign xor_ln28_20_fu_4982_p2 = (z2_50_fu_4956_p2 ^ z1_52_fu_4950_p2);

assign xor_ln28_21_fu_5040_p2 = (a1_92_fu_5032_p3 ^ a0_105_fu_5028_p1);

assign xor_ln28_22_fu_5054_p2 = (tmp_20_fu_5046_p3 ^ a0_103_fu_5014_p2);

assign xor_ln28_23_fu_5514_p2 = (z2_55_fu_5488_p2 ^ z1_56_fu_5482_p2);

assign xor_ln28_24_fu_5890_p2 = (z2_59_fu_5864_p2 ^ z1_60_fu_5858_p2);

assign xor_ln28_25_fu_6194_p2 = (z2_63_fu_6168_p2 ^ z1_65_fu_6162_p2);

assign xor_ln28_26_fu_6252_p2 = (a1_114_fu_6244_p3 ^ a0_131_fu_6240_p1);

assign xor_ln28_27_fu_6266_p2 = (tmp_25_fu_6258_p3 ^ a0_130_fu_6226_p2);

assign xor_ln28_28_fu_6590_p2 = (z2_68_fu_6564_p2 ^ z1_70_fu_6558_p2);

assign xor_ln28_29_fu_6966_p2 = (z2_72_fu_6940_p2 ^ z1_74_fu_6934_p2);

assign xor_ln28_2_fu_1230_p2 = (z2_10_fu_1204_p2 ^ z1_12_fu_1198_p2);

assign xor_ln28_30_fu_7270_p2 = (z2_76_fu_7244_p2 ^ z1_79_fu_7238_p2);

assign xor_ln28_31_fu_7328_p2 = (a1_135_fu_7320_p3 ^ a0_146_fu_7316_p1);

assign xor_ln28_32_fu_7342_p2 = (tmp_30_fu_7334_p3 ^ a0_145_fu_7302_p2);

assign xor_ln28_33_fu_7418_p2 = (a1_138_fu_7410_p3 ^ a0_149_fu_7402_p3);

assign xor_ln28_34_fu_7432_p2 = (tmp_32_fu_7424_p3 ^ a0_148_fu_7388_p1);

assign xor_ln28_35_fu_7446_p2 = (tmp_33_fu_7438_p3 ^ a0_147_fu_7374_p2);

assign xor_ln28_36_fu_7790_p2 = (z2_82_fu_7764_p2 ^ z1_84_fu_7758_p2);

assign xor_ln28_37_fu_8166_p2 = (z2_86_fu_8140_p2 ^ z1_88_fu_8134_p2);

assign xor_ln28_38_fu_8470_p2 = (z2_90_fu_8444_p2 ^ z1_93_fu_8438_p2);

assign xor_ln28_39_fu_8528_p2 = (a1_161_fu_8520_p3 ^ a0_166_fu_8516_p1);

assign xor_ln28_3_fu_1288_p2 = (a1_23_fu_1280_p3 ^ a0_23_fu_1276_p1);

assign xor_ln28_40_fu_8542_p2 = (tmp_38_fu_8534_p3 ^ a0_165_fu_8502_p2);

assign xor_ln28_41_fu_9002_p2 = (z2_95_fu_8976_p2 ^ z1_97_fu_8970_p2);

assign xor_ln28_42_fu_9378_p2 = (z2_99_fu_9352_p2 ^ z1_101_fu_9346_p2);

assign xor_ln28_43_fu_9682_p2 = (z2_103_fu_9656_p2 ^ z1_106_fu_9650_p2);

assign xor_ln28_44_fu_9740_p2 = (a1_180_fu_9732_p3 ^ a0_183_fu_9728_p1);

assign xor_ln28_45_fu_9754_p2 = (tmp_43_fu_9746_p3 ^ a0_182_fu_9714_p2);

assign xor_ln28_46_fu_10078_p2 = (z2_108_fu_10052_p2 ^ z1_111_fu_10046_p2);

assign xor_ln28_47_fu_10454_p2 = (z2_112_fu_10428_p2 ^ z1_115_fu_10422_p2);

assign xor_ln28_48_fu_10758_p2 = (z2_116_fu_10732_p2 ^ z1_120_fu_10726_p2);

assign xor_ln28_49_fu_10816_p2 = (a1_197_fu_10808_p3 ^ a0_200_fu_10804_p1);

assign xor_ln28_4_fu_1302_p2 = (tmp_1_fu_1294_p3 ^ a0_21_fu_1262_p2);

assign xor_ln28_50_fu_10830_p2 = (tmp_48_fu_10822_p3 ^ a0_199_fu_10790_p2);

assign xor_ln28_51_fu_10906_p2 = (a1_200_fu_10898_p3 ^ a0_203_fu_10890_p3);

assign xor_ln28_52_fu_10920_p2 = (tmp_50_fu_10912_p3 ^ a0_202_fu_10876_p1);

assign xor_ln28_53_fu_10934_p2 = (tmp_51_fu_10926_p3 ^ a0_201_fu_10862_p2);

assign xor_ln28_54_fu_11030_p2 = (a1_204_fu_11022_p3 ^ a0_207_fu_11014_p3);

assign xor_ln28_55_fu_11044_p2 = (tmp_53_fu_11036_p3 ^ a0_206_fu_10994_p4);

assign xor_ln28_56_fu_11058_p2 = (tmp_54_fu_11050_p3 ^ a0_205_fu_10980_p1);

assign xor_ln28_57_fu_11072_p2 = (tmp_55_fu_11064_p3 ^ a0_204_fu_10966_p2);

assign xor_ln28_5_fu_1762_p2 = (z2_15_fu_1736_p2 ^ z1_16_fu_1730_p2);

assign xor_ln28_6_fu_2138_p2 = (z2_19_fu_2112_p2 ^ z1_20_fu_2106_p2);

assign xor_ln28_7_fu_2442_p2 = (z2_23_fu_2416_p2 ^ z1_25_fu_2410_p2);

assign xor_ln28_8_fu_2500_p2 = (a1_45_fu_2492_p3 ^ a0_48_fu_2488_p1);

assign xor_ln28_9_fu_2514_p2 = (tmp_7_fu_2506_p3 ^ a0_47_fu_2474_p2);

assign xor_ln28_fu_550_p2 = (z2_2_fu_524_p2 ^ z1_3_fu_518_p2);

assign xor_ln33_1_fu_3906_p2 = (trunc_ln43_7_fu_3890_p4 ^ trunc_ln40_1_fu_190_p1);

assign xor_ln33_2_fu_3912_p2 = (trunc_ln43_6_fu_3880_p4 ^ trunc_ln40_2_fu_194_p1);

assign xor_ln33_3_fu_3918_p2 = (trunc_ln43_5_fu_3870_p4 ^ trunc_ln40_3_fu_198_p1);

assign xor_ln33_4_fu_5194_p2 = (xor_ln40_1_fu_3972_p2 ^ trunc_ln43_9_fu_5178_p4);

assign xor_ln33_5_fu_8682_p2 = (trunc_ln43_11_fu_8666_p4 ^ trunc_ln40_5_fu_3956_p4);

assign xor_ln33_fu_1442_p2 = (trunc_ln43_1_fu_1426_p4 ^ trunc_ln40_4_fu_234_p1);

assign xor_ln38_1_fu_3940_p2 = (trunc_ln38_5_fu_3924_p4 ^ trunc_ln38_4_fu_216_p1);

assign xor_ln40_1_fu_3972_p2 = (trunc_ln40_5_fu_3956_p4 ^ trunc_ln40_4_fu_234_p1);

assign xor_ln43_100_fu_8632_p2 = (trunc_ln43_10_fu_8616_p4 ^ trunc_ln38_5_fu_3924_p4);

assign xor_ln43_14_fu_1392_p2 = (trunc_ln43_s_fu_1376_p4 ^ trunc_ln38_4_fu_216_p1);

assign xor_ln43_42_fu_3814_p2 = (trunc_ln43_4_fu_3798_p4 ^ trunc_ln38_1_fu_164_p1);

assign xor_ln43_43_fu_3820_p2 = (trunc_ln43_3_fu_3788_p4 ^ trunc_ln38_2_fu_168_p1);

assign xor_ln43_44_fu_3826_p2 = (trunc_ln43_2_fu_3778_p4 ^ trunc_ln38_3_fu_172_p1);

assign xor_ln43_59_fu_5144_p2 = (xor_ln38_1_fu_3940_p2 ^ trunc_ln43_8_fu_5128_p4);

assign xor_ln45_102_fu_3708_p2 = (z1_26_fu_2552_p3 ^ z0_13_fu_1340_p3);

assign xor_ln45_103_fu_3714_p2 = (z2_133_fu_3628_p3 ^ tmp_16_fu_3700_p3);

assign xor_ln45_104_fu_3720_p2 = (xor_ln45_103_fu_3714_p2 ^ xor_ln45_102_fu_3708_p2);

assign xor_ln45_105_fu_3726_p2 = (z2_133_fu_3628_p3 ^ z0_13_fu_1340_p3);

assign xor_ln45_106_fu_4110_p2 = (z1_40_fu_4098_p2 ^ z0_41_fu_4080_p2);

assign xor_ln45_107_fu_4116_p2 = (z2_40_fu_4104_p2 ^ z0_41_fu_4080_p2);

assign xor_ln45_108_fu_4216_p2 = (z1_41_fu_4204_p2 ^ z0_43_fu_4186_p2);

assign xor_ln45_109_fu_4222_p2 = (z2_41_fu_4210_p2 ^ z0_43_fu_4186_p2);

assign xor_ln45_10_fu_734_p2 = (z1_4_fu_722_p2 ^ z0_5_fu_704_p2);

assign xor_ln45_112_fu_4316_p2 = (z1_42_fu_4228_p3 ^ z0_42_fu_4122_p3);

assign xor_ln45_113_fu_4322_p2 = (z2_134_fu_4294_p3 ^ tmp_17_fu_4308_p3);

assign xor_ln45_114_fu_4328_p2 = (xor_ln45_113_fu_4322_p2 ^ xor_ln45_112_fu_4316_p2);

assign xor_ln45_115_fu_4334_p2 = (z2_134_fu_4294_p3 ^ z0_42_fu_4122_p3);

assign xor_ln45_116_fu_4486_p2 = (z1_44_fu_4474_p2 ^ z0_46_fu_4456_p2);

assign xor_ln45_117_fu_4492_p2 = (z2_44_fu_4480_p2 ^ z0_46_fu_4456_p2);

assign xor_ln45_118_fu_4592_p2 = (z1_45_fu_4580_p2 ^ z0_48_fu_4562_p2);

assign xor_ln45_119_fu_4598_p2 = (z2_45_fu_4586_p2 ^ z0_48_fu_4562_p2);

assign xor_ln45_11_fu_740_p2 = (z2_4_fu_728_p2 ^ z0_5_fu_704_p2);

assign xor_ln45_122_fu_4692_p2 = (z1_46_fu_4604_p3 ^ z0_47_fu_4498_p3);

assign xor_ln45_123_fu_4698_p2 = (z2_135_fu_4670_p3 ^ tmp_18_fu_4684_p3);

assign xor_ln45_124_fu_4704_p2 = (xor_ln45_123_fu_4698_p2 ^ xor_ln45_122_fu_4692_p2);

assign xor_ln45_125_fu_4710_p2 = (z2_135_fu_4670_p3 ^ z0_47_fu_4498_p3);

assign xor_ln45_126_fu_4790_p2 = (z1_49_fu_4778_p2 ^ z0_50_fu_4760_p2);

assign xor_ln45_127_fu_4796_p2 = (z2_48_fu_4784_p2 ^ z0_50_fu_4760_p2);

assign xor_ln45_128_fu_4896_p2 = (z1_50_fu_4884_p2 ^ z0_52_fu_4866_p2);

assign xor_ln45_129_fu_4902_p2 = (z2_49_fu_4890_p2 ^ z0_52_fu_4866_p2);

assign xor_ln45_12_fu_840_p2 = (z1_5_fu_828_p2 ^ z0_7_fu_810_p2);

assign xor_ln45_132_fu_4996_p2 = (z1_51_fu_4908_p3 ^ z0_51_fu_4802_p3);

assign xor_ln45_133_fu_5002_p2 = (z2_136_fu_4974_p3 ^ tmp_19_fu_4988_p3);

assign xor_ln45_136_fu_5068_p2 = (z1_48_fu_4716_p3 ^ z0_45_fu_4340_p3);

assign xor_ln45_137_fu_5074_p2 = (z2_137_fu_5020_p3 ^ tmp_21_fu_5060_p3);

assign xor_ln45_138_fu_5080_p2 = (xor_ln45_137_fu_5074_p2 ^ xor_ln45_136_fu_5068_p2);

assign xor_ln45_139_fu_5086_p2 = (z2_137_fu_5020_p3 ^ z0_45_fu_4340_p3);

assign xor_ln45_13_fu_846_p2 = (z2_5_fu_834_p2 ^ z0_7_fu_810_p2);

assign xor_ln45_140_fu_5322_p2 = (z1_53_fu_5310_p2 ^ z0_55_fu_5292_p2);

assign xor_ln45_141_fu_5328_p2 = (z2_53_fu_5316_p2 ^ z0_55_fu_5292_p2);

assign xor_ln45_142_fu_5428_p2 = (z1_54_fu_5416_p2 ^ z0_57_fu_5398_p2);

assign xor_ln45_143_fu_5434_p2 = (z2_54_fu_5422_p2 ^ z0_57_fu_5398_p2);

assign xor_ln45_146_fu_5528_p2 = (z1_55_fu_5440_p3 ^ z0_56_fu_5334_p3);

assign xor_ln45_147_fu_5534_p2 = (z2_138_fu_5506_p3 ^ tmp_22_fu_5520_p3);

assign xor_ln45_148_fu_5540_p2 = (xor_ln45_147_fu_5534_p2 ^ xor_ln45_146_fu_5528_p2);

assign xor_ln45_149_fu_5546_p2 = (z2_138_fu_5506_p3 ^ z0_56_fu_5334_p3);

assign xor_ln45_150_fu_5698_p2 = (z1_57_fu_5686_p2 ^ z0_60_fu_5668_p2);

assign xor_ln45_151_fu_5704_p2 = (z2_57_fu_5692_p2 ^ z0_60_fu_5668_p2);

assign xor_ln45_152_fu_5804_p2 = (z1_58_fu_5792_p2 ^ z0_62_fu_5774_p2);

assign xor_ln45_153_fu_5810_p2 = (z2_58_fu_5798_p2 ^ z0_62_fu_5774_p2);

assign xor_ln45_156_fu_5904_p2 = (z1_59_fu_5816_p3 ^ z0_61_fu_5710_p3);

assign xor_ln45_157_fu_5910_p2 = (z2_139_fu_5882_p3 ^ tmp_23_fu_5896_p3);

assign xor_ln45_158_fu_5916_p2 = (xor_ln45_157_fu_5910_p2 ^ xor_ln45_156_fu_5904_p2);

assign xor_ln45_159_fu_5922_p2 = (z2_139_fu_5882_p3 ^ z0_61_fu_5710_p3);

assign xor_ln45_160_fu_6002_p2 = (z1_62_fu_5990_p2 ^ z0_64_fu_5972_p2);

assign xor_ln45_161_fu_6008_p2 = (z2_61_fu_5996_p2 ^ z0_64_fu_5972_p2);

assign xor_ln45_162_fu_6108_p2 = (z1_63_fu_6096_p2 ^ z0_66_fu_6078_p2);

assign xor_ln45_163_fu_6114_p2 = (z2_62_fu_6102_p2 ^ z0_66_fu_6078_p2);

assign xor_ln45_166_fu_6208_p2 = (z1_64_fu_6120_p3 ^ z0_65_fu_6014_p3);

assign xor_ln45_167_fu_6214_p2 = (z2_140_fu_6186_p3 ^ tmp_24_fu_6200_p3);

assign xor_ln45_16_fu_940_p2 = (z1_6_fu_852_p3 ^ z0_6_fu_746_p3);

assign xor_ln45_170_fu_6280_p2 = (z1_61_fu_5928_p3 ^ z0_59_fu_5552_p3);

assign xor_ln45_171_fu_6286_p2 = (z2_141_fu_6232_p3 ^ tmp_26_fu_6272_p3);

assign xor_ln45_172_fu_6292_p2 = (xor_ln45_171_fu_6286_p2 ^ xor_ln45_170_fu_6280_p2);

assign xor_ln45_173_fu_6298_p2 = (z2_141_fu_6232_p3 ^ z0_59_fu_5552_p3);

assign xor_ln45_174_fu_6398_p2 = (z1_67_fu_6386_p2 ^ z0_68_fu_6368_p2);

assign xor_ln45_175_fu_6404_p2 = (z2_66_fu_6392_p2 ^ z0_68_fu_6368_p2);

assign xor_ln45_176_fu_6504_p2 = (z1_68_fu_6492_p2 ^ z0_70_fu_6474_p2);

assign xor_ln45_177_fu_6510_p2 = (z2_67_fu_6498_p2 ^ z0_70_fu_6474_p2);

assign xor_ln45_17_fu_946_p2 = (z2_122_fu_918_p3 ^ tmp_5_fu_932_p3);

assign xor_ln45_180_fu_6604_p2 = (z1_69_fu_6516_p3 ^ z0_69_fu_6410_p3);

assign xor_ln45_181_fu_6610_p2 = (z2_142_fu_6582_p3 ^ tmp_27_fu_6596_p3);

assign xor_ln45_182_fu_6616_p2 = (xor_ln45_181_fu_6610_p2 ^ xor_ln45_180_fu_6604_p2);

assign xor_ln45_183_fu_6622_p2 = (z2_142_fu_6582_p3 ^ z0_69_fu_6410_p3);

assign xor_ln45_184_fu_6774_p2 = (z1_71_fu_6762_p2 ^ z0_73_fu_6744_p2);

assign xor_ln45_185_fu_6780_p2 = (z2_70_fu_6768_p2 ^ z0_73_fu_6744_p2);

assign xor_ln45_186_fu_6880_p2 = (z1_72_fu_6868_p2 ^ z0_75_fu_6850_p2);

assign xor_ln45_187_fu_6886_p2 = (z2_71_fu_6874_p2 ^ z0_75_fu_6850_p2);

assign xor_ln45_18_fu_952_p2 = (xor_ln45_17_fu_946_p2 ^ xor_ln45_16_fu_940_p2);

assign xor_ln45_190_fu_6980_p2 = (z1_73_fu_6892_p3 ^ z0_74_fu_6786_p3);

assign xor_ln45_191_fu_6986_p2 = (z2_143_fu_6958_p3 ^ tmp_28_fu_6972_p3);

assign xor_ln45_192_fu_6992_p2 = (xor_ln45_191_fu_6986_p2 ^ xor_ln45_190_fu_6980_p2);

assign xor_ln45_193_fu_6998_p2 = (z2_143_fu_6958_p3 ^ z0_74_fu_6786_p3);

assign xor_ln45_194_fu_7078_p2 = (z1_76_fu_7066_p2 ^ z0_77_fu_7048_p2);

assign xor_ln45_195_fu_7084_p2 = (z2_74_fu_7072_p2 ^ z0_77_fu_7048_p2);

assign xor_ln45_196_fu_7184_p2 = (z1_77_fu_7172_p2 ^ z0_79_fu_7154_p2);

assign xor_ln45_197_fu_7190_p2 = (z2_75_fu_7178_p2 ^ z0_79_fu_7154_p2);

assign xor_ln45_19_fu_958_p2 = (z2_122_fu_918_p3 ^ z0_6_fu_746_p3);

assign xor_ln45_1_fu_364_p2 = (z2_fu_352_p2 ^ z0_fu_328_p2);

assign xor_ln45_200_fu_7284_p2 = (z1_78_fu_7196_p3 ^ z0_78_fu_7090_p3);

assign xor_ln45_201_fu_7290_p2 = (z2_144_fu_7262_p3 ^ tmp_29_fu_7276_p3);

assign xor_ln45_204_fu_7356_p2 = (z1_75_fu_7004_p3 ^ z0_72_fu_6628_p3);

assign xor_ln45_205_fu_7362_p2 = (z2_145_fu_7308_p3 ^ tmp_31_fu_7348_p3);

assign xor_ln45_208_fu_7460_p2 = (z1_66_fu_6304_p3 ^ z0_54_fu_5092_p3);

assign xor_ln45_209_fu_7466_p2 = (z2_146_fu_7380_p3 ^ tmp_34_fu_7452_p3);

assign xor_ln45_20_fu_1038_p2 = (z1_9_fu_1026_p2 ^ z0_9_fu_1008_p2);

assign xor_ln45_210_fu_7472_p2 = (xor_ln45_209_fu_7466_p2 ^ xor_ln45_208_fu_7460_p2);

assign xor_ln45_211_fu_7478_p2 = (z2_146_fu_7380_p3 ^ z0_54_fu_5092_p3);

assign xor_ln45_212_fu_7598_p2 = (z1_81_fu_7586_p2 ^ z0_81_fu_7568_p2);

assign xor_ln45_213_fu_7604_p2 = (z2_80_fu_7592_p2 ^ z0_81_fu_7568_p2);

assign xor_ln45_214_fu_7704_p2 = (z1_82_fu_7692_p2 ^ z0_83_fu_7674_p2);

assign xor_ln45_215_fu_7710_p2 = (z2_81_fu_7698_p2 ^ z0_83_fu_7674_p2);

assign xor_ln45_218_fu_7804_p2 = (z1_83_fu_7716_p3 ^ z0_82_fu_7610_p3);

assign xor_ln45_219_fu_7810_p2 = (z2_147_fu_7782_p3 ^ tmp_35_fu_7796_p3);

assign xor_ln45_21_fu_1044_p2 = (z2_8_fu_1032_p2 ^ z0_9_fu_1008_p2);

assign xor_ln45_220_fu_7816_p2 = (xor_ln45_219_fu_7810_p2 ^ xor_ln45_218_fu_7804_p2);

assign xor_ln45_221_fu_7822_p2 = (z2_147_fu_7782_p3 ^ z0_82_fu_7610_p3);

assign xor_ln45_222_fu_7974_p2 = (z1_85_fu_7962_p2 ^ z0_86_fu_7944_p2);

assign xor_ln45_223_fu_7980_p2 = (z2_84_fu_7968_p2 ^ z0_86_fu_7944_p2);

assign xor_ln45_224_fu_8080_p2 = (z1_86_fu_8068_p2 ^ z0_88_fu_8050_p2);

assign xor_ln45_225_fu_8086_p2 = (z2_85_fu_8074_p2 ^ z0_88_fu_8050_p2);

assign xor_ln45_228_fu_8180_p2 = (z1_87_fu_8092_p3 ^ z0_87_fu_7986_p3);

assign xor_ln45_229_fu_8186_p2 = (z2_148_fu_8158_p3 ^ tmp_36_fu_8172_p3);

assign xor_ln45_22_fu_1144_p2 = (z1_10_fu_1132_p2 ^ z0_11_fu_1114_p2);

assign xor_ln45_230_fu_8192_p2 = (xor_ln45_229_fu_8186_p2 ^ xor_ln45_228_fu_8180_p2);

assign xor_ln45_231_fu_8198_p2 = (z2_148_fu_8158_p3 ^ z0_87_fu_7986_p3);

assign xor_ln45_232_fu_8278_p2 = (z1_90_fu_8266_p2 ^ z0_90_fu_8248_p2);

assign xor_ln45_233_fu_8284_p2 = (z2_88_fu_8272_p2 ^ z0_90_fu_8248_p2);

assign xor_ln45_234_fu_8384_p2 = (z1_91_fu_8372_p2 ^ z0_92_fu_8354_p2);

assign xor_ln45_235_fu_8390_p2 = (z2_89_fu_8378_p2 ^ z0_92_fu_8354_p2);

assign xor_ln45_238_fu_8484_p2 = (z1_92_fu_8396_p3 ^ z0_91_fu_8290_p3);

assign xor_ln45_239_fu_8490_p2 = (z2_149_fu_8462_p3 ^ tmp_37_fu_8476_p3);

assign xor_ln45_23_fu_1150_p2 = (z2_9_fu_1138_p2 ^ z0_11_fu_1114_p2);

assign xor_ln45_242_fu_8556_p2 = (z1_89_fu_8204_p3 ^ z0_85_fu_7828_p3);

assign xor_ln45_243_fu_8562_p2 = (z2_150_fu_8508_p3 ^ tmp_39_fu_8548_p3);

assign xor_ln45_244_fu_8568_p2 = (xor_ln45_243_fu_8562_p2 ^ xor_ln45_242_fu_8556_p2);

assign xor_ln45_245_fu_8574_p2 = (z2_150_fu_8508_p3 ^ z0_85_fu_7828_p3);

assign xor_ln45_246_fu_8810_p2 = (z1_94_fu_8798_p2 ^ z0_95_fu_8780_p2);

assign xor_ln45_247_fu_8816_p2 = (z2_93_fu_8804_p2 ^ z0_95_fu_8780_p2);

assign xor_ln45_248_fu_8916_p2 = (z1_95_fu_8904_p2 ^ z0_97_fu_8886_p2);

assign xor_ln45_249_fu_8922_p2 = (z2_94_fu_8910_p2 ^ z0_97_fu_8886_p2);

assign xor_ln45_252_fu_9016_p2 = (z1_96_fu_8928_p3 ^ z0_96_fu_8822_p3);

assign xor_ln45_253_fu_9022_p2 = (z2_151_fu_8994_p3 ^ tmp_40_fu_9008_p3);

assign xor_ln45_254_fu_9028_p2 = (xor_ln45_253_fu_9022_p2 ^ xor_ln45_252_fu_9016_p2);

assign xor_ln45_255_fu_9034_p2 = (z2_151_fu_8994_p3 ^ z0_96_fu_8822_p3);

assign xor_ln45_256_fu_9186_p2 = (z1_98_fu_9174_p2 ^ z0_100_fu_9156_p2);

assign xor_ln45_257_fu_9192_p2 = (z2_97_fu_9180_p2 ^ z0_100_fu_9156_p2);

assign xor_ln45_258_fu_9292_p2 = (z1_99_fu_9280_p2 ^ z0_102_fu_9262_p2);

assign xor_ln45_259_fu_9298_p2 = (z2_98_fu_9286_p2 ^ z0_102_fu_9262_p2);

assign xor_ln45_262_fu_9392_p2 = (z1_100_fu_9304_p3 ^ z0_101_fu_9198_p3);

assign xor_ln45_263_fu_9398_p2 = (z2_152_fu_9370_p3 ^ tmp_41_fu_9384_p3);

assign xor_ln45_264_fu_9404_p2 = (xor_ln45_263_fu_9398_p2 ^ xor_ln45_262_fu_9392_p2);

assign xor_ln45_265_fu_9410_p2 = (z2_152_fu_9370_p3 ^ z0_101_fu_9198_p3);

assign xor_ln45_266_fu_9490_p2 = (z1_103_fu_9478_p2 ^ z0_104_fu_9460_p2);

assign xor_ln45_267_fu_9496_p2 = (z2_101_fu_9484_p2 ^ z0_104_fu_9460_p2);

assign xor_ln45_268_fu_9596_p2 = (z1_104_fu_9584_p2 ^ z0_106_fu_9566_p2);

assign xor_ln45_269_fu_9602_p2 = (z2_102_fu_9590_p2 ^ z0_106_fu_9566_p2);

assign xor_ln45_26_fu_1244_p2 = (z1_11_fu_1156_p3 ^ z0_10_fu_1050_p3);

assign xor_ln45_272_fu_9696_p2 = (z1_105_fu_9608_p3 ^ z0_105_fu_9502_p3);

assign xor_ln45_273_fu_9702_p2 = (z2_153_fu_9674_p3 ^ tmp_42_fu_9688_p3);

assign xor_ln45_276_fu_9768_p2 = (z1_102_fu_9416_p3 ^ z0_99_fu_9040_p3);

assign xor_ln45_277_fu_9774_p2 = (z2_154_fu_9720_p3 ^ tmp_44_fu_9760_p3);

assign xor_ln45_278_fu_9780_p2 = (xor_ln45_277_fu_9774_p2 ^ xor_ln45_276_fu_9768_p2);

assign xor_ln45_279_fu_9786_p2 = (z2_154_fu_9720_p3 ^ z0_99_fu_9040_p3);

assign xor_ln45_27_fu_1250_p2 = (z2_123_fu_1222_p3 ^ tmp_s_fu_1236_p3);

assign xor_ln45_280_fu_9886_p2 = (z1_108_fu_9874_p2 ^ z0_108_fu_9856_p2);

assign xor_ln45_281_fu_9892_p2 = (z2_106_fu_9880_p2 ^ z0_108_fu_9856_p2);

assign xor_ln45_282_fu_9992_p2 = (z1_109_fu_9980_p2 ^ z0_110_fu_9962_p2);

assign xor_ln45_283_fu_9998_p2 = (z2_107_fu_9986_p2 ^ z0_110_fu_9962_p2);

assign xor_ln45_286_fu_10092_p2 = (z1_110_fu_10004_p3 ^ z0_109_fu_9898_p3);

assign xor_ln45_287_fu_10098_p2 = (z2_155_fu_10070_p3 ^ tmp_45_fu_10084_p3);

assign xor_ln45_288_fu_10104_p2 = (xor_ln45_287_fu_10098_p2 ^ xor_ln45_286_fu_10092_p2);

assign xor_ln45_289_fu_10110_p2 = (z2_155_fu_10070_p3 ^ z0_109_fu_9898_p3);

assign xor_ln45_290_fu_10262_p2 = (z1_112_fu_10250_p2 ^ z0_113_fu_10232_p2);

assign xor_ln45_291_fu_10268_p2 = (z2_110_fu_10256_p2 ^ z0_113_fu_10232_p2);

assign xor_ln45_292_fu_10368_p2 = (z1_113_fu_10356_p2 ^ z0_115_fu_10338_p2);

assign xor_ln45_293_fu_10374_p2 = (z2_111_fu_10362_p2 ^ z0_115_fu_10338_p2);

assign xor_ln45_296_fu_10468_p2 = (z1_114_fu_10380_p3 ^ z0_114_fu_10274_p3);

assign xor_ln45_297_fu_10474_p2 = (z2_156_fu_10446_p3 ^ tmp_46_fu_10460_p3);

assign xor_ln45_298_fu_10480_p2 = (xor_ln45_297_fu_10474_p2 ^ xor_ln45_296_fu_10468_p2);

assign xor_ln45_299_fu_10486_p2 = (z2_156_fu_10446_p3 ^ z0_114_fu_10274_p3);

assign xor_ln45_2_fu_464_p2 = (z1_1_fu_452_p2 ^ z0_2_fu_434_p2);

assign xor_ln45_300_fu_10566_p2 = (z1_117_fu_10554_p2 ^ z0_117_fu_10536_p2);

assign xor_ln45_301_fu_10572_p2 = (z2_114_fu_10560_p2 ^ z0_117_fu_10536_p2);

assign xor_ln45_302_fu_10672_p2 = (z1_118_fu_10660_p2 ^ z0_119_fu_10642_p2);

assign xor_ln45_303_fu_10678_p2 = (z2_115_fu_10666_p2 ^ z0_119_fu_10642_p2);

assign xor_ln45_306_fu_10772_p2 = (z1_119_fu_10684_p3 ^ z0_118_fu_10578_p3);

assign xor_ln45_307_fu_10778_p2 = (z2_157_fu_10750_p3 ^ tmp_47_fu_10764_p3);

assign xor_ln45_30_fu_1316_p2 = (z1_8_fu_964_p3 ^ z0_4_fu_588_p3);

assign xor_ln45_310_fu_10844_p2 = (z1_116_fu_10492_p3 ^ z0_112_fu_10116_p3);

assign xor_ln45_311_fu_10850_p2 = (z2_158_fu_10796_p3 ^ tmp_49_fu_10836_p3);

assign xor_ln45_314_fu_10948_p2 = (z1_107_fu_9792_p3 ^ z0_94_fu_8580_p3);

assign xor_ln45_315_fu_10954_p2 = (z2_159_fu_10868_p3 ^ tmp_52_fu_10940_p3);

assign xor_ln45_318_fu_11086_p2 = (z1_80_fu_7484_p3 ^ z0_40_fu_3732_p3);

assign xor_ln45_319_fu_11092_p2 = (z2_160_fu_10972_p3 ^ tmp_56_fu_11078_p3);

assign xor_ln45_31_fu_1322_p2 = (z2_124_fu_1268_p3 ^ tmp_2_fu_1308_p3);

assign xor_ln45_320_fu_11098_p2 = (xor_ln45_319_fu_11092_p2 ^ xor_ln45_318_fu_11086_p2);

assign xor_ln45_321_fu_11104_p2 = (z2_160_fu_10972_p3 ^ z0_40_fu_3732_p3);

assign xor_ln45_32_fu_1328_p2 = (xor_ln45_31_fu_1322_p2 ^ xor_ln45_30_fu_1316_p2);

assign xor_ln45_33_fu_1334_p2 = (z2_124_fu_1268_p3 ^ z0_4_fu_588_p3);

assign xor_ln45_34_fu_1570_p2 = (z1_13_fu_1558_p2 ^ z0_14_fu_1540_p2);

assign xor_ln45_35_fu_1576_p2 = (z2_13_fu_1564_p2 ^ z0_14_fu_1540_p2);

assign xor_ln45_36_fu_1676_p2 = (z1_14_fu_1664_p2 ^ z0_16_fu_1646_p2);

assign xor_ln45_37_fu_1682_p2 = (z2_14_fu_1670_p2 ^ z0_16_fu_1646_p2);

assign xor_ln45_3_fu_470_p2 = (z2_1_fu_458_p2 ^ z0_2_fu_434_p2);

assign xor_ln45_40_fu_1776_p2 = (z1_15_fu_1688_p3 ^ z0_15_fu_1582_p3);

assign xor_ln45_41_fu_1782_p2 = (z2_125_fu_1754_p3 ^ tmp_3_fu_1768_p3);

assign xor_ln45_42_fu_1788_p2 = (xor_ln45_41_fu_1782_p2 ^ xor_ln45_40_fu_1776_p2);

assign xor_ln45_43_fu_1794_p2 = (z2_125_fu_1754_p3 ^ z0_15_fu_1582_p3);

assign xor_ln45_44_fu_1946_p2 = (z1_17_fu_1934_p2 ^ z0_19_fu_1916_p2);

assign xor_ln45_45_fu_1952_p2 = (z2_17_fu_1940_p2 ^ z0_19_fu_1916_p2);

assign xor_ln45_46_fu_2052_p2 = (z1_18_fu_2040_p2 ^ z0_21_fu_2022_p2);

assign xor_ln45_47_fu_2058_p2 = (z2_18_fu_2046_p2 ^ z0_21_fu_2022_p2);

assign xor_ln45_50_fu_2152_p2 = (z1_19_fu_2064_p3 ^ z0_20_fu_1958_p3);

assign xor_ln45_51_fu_2158_p2 = (z2_126_fu_2130_p3 ^ tmp_4_fu_2144_p3);

assign xor_ln45_52_fu_2164_p2 = (xor_ln45_51_fu_2158_p2 ^ xor_ln45_50_fu_2152_p2);

assign xor_ln45_53_fu_2170_p2 = (z2_126_fu_2130_p3 ^ z0_20_fu_1958_p3);

assign xor_ln45_54_fu_2250_p2 = (z1_22_fu_2238_p2 ^ z0_23_fu_2220_p2);

assign xor_ln45_55_fu_2256_p2 = (z2_21_fu_2244_p2 ^ z0_23_fu_2220_p2);

assign xor_ln45_56_fu_2356_p2 = (z1_23_fu_2344_p2 ^ z0_25_fu_2326_p2);

assign xor_ln45_57_fu_2362_p2 = (z2_22_fu_2350_p2 ^ z0_25_fu_2326_p2);

assign xor_ln45_60_fu_2456_p2 = (z1_24_fu_2368_p3 ^ z0_24_fu_2262_p3);

assign xor_ln45_61_fu_2462_p2 = (z2_127_fu_2434_p3 ^ tmp_6_fu_2448_p3);

assign xor_ln45_64_fu_2528_p2 = (z1_21_fu_2176_p3 ^ z0_18_fu_1800_p3);

assign xor_ln45_65_fu_2534_p2 = (z2_128_fu_2480_p3 ^ tmp_8_fu_2520_p3);

assign xor_ln45_66_fu_2540_p2 = (xor_ln45_65_fu_2534_p2 ^ xor_ln45_64_fu_2528_p2);

assign xor_ln45_67_fu_2546_p2 = (z2_128_fu_2480_p3 ^ z0_18_fu_1800_p3);

assign xor_ln45_68_fu_2646_p2 = (z1_27_fu_2634_p2 ^ z0_27_fu_2616_p2);

assign xor_ln45_69_fu_2652_p2 = (z2_26_fu_2640_p2 ^ z0_27_fu_2616_p2);

assign xor_ln45_6_fu_564_p2 = (z1_2_fu_476_p3 ^ z0_1_fu_370_p3);

assign xor_ln45_70_fu_2752_p2 = (z1_28_fu_2740_p2 ^ z0_29_fu_2722_p2);

assign xor_ln45_71_fu_2758_p2 = (z2_27_fu_2746_p2 ^ z0_29_fu_2722_p2);

assign xor_ln45_74_fu_2852_p2 = (z1_29_fu_2764_p3 ^ z0_28_fu_2658_p3);

assign xor_ln45_75_fu_2858_p2 = (z2_129_fu_2830_p3 ^ tmp_9_fu_2844_p3);

assign xor_ln45_76_fu_2864_p2 = (xor_ln45_75_fu_2858_p2 ^ xor_ln45_74_fu_2852_p2);

assign xor_ln45_77_fu_2870_p2 = (z2_129_fu_2830_p3 ^ z0_28_fu_2658_p3);

assign xor_ln45_78_fu_3022_p2 = (z1_31_fu_3010_p2 ^ z0_32_fu_2992_p2);

assign xor_ln45_79_fu_3028_p2 = (z2_30_fu_3016_p2 ^ z0_32_fu_2992_p2);

assign xor_ln45_7_fu_570_p2 = (z2_121_fu_542_p3 ^ tmp_fu_556_p3);

assign xor_ln45_80_fu_3128_p2 = (z1_32_fu_3116_p2 ^ z0_34_fu_3098_p2);

assign xor_ln45_81_fu_3134_p2 = (z2_31_fu_3122_p2 ^ z0_34_fu_3098_p2);

assign xor_ln45_84_fu_3228_p2 = (z1_33_fu_3140_p3 ^ z0_33_fu_3034_p3);

assign xor_ln45_85_fu_3234_p2 = (z2_130_fu_3206_p3 ^ tmp_10_fu_3220_p3);

assign xor_ln45_86_fu_3240_p2 = (xor_ln45_85_fu_3234_p2 ^ xor_ln45_84_fu_3228_p2);

assign xor_ln45_87_fu_3246_p2 = (z2_130_fu_3206_p3 ^ z0_33_fu_3034_p3);

assign xor_ln45_88_fu_3326_p2 = (z1_36_fu_3314_p2 ^ z0_36_fu_3296_p2);

assign xor_ln45_89_fu_3332_p2 = (z2_34_fu_3320_p2 ^ z0_36_fu_3296_p2);

assign xor_ln45_8_fu_576_p2 = (xor_ln45_7_fu_570_p2 ^ xor_ln45_6_fu_564_p2);

assign xor_ln45_90_fu_3432_p2 = (z1_37_fu_3420_p2 ^ z0_38_fu_3402_p2);

assign xor_ln45_91_fu_3438_p2 = (z2_35_fu_3426_p2 ^ z0_38_fu_3402_p2);

assign xor_ln45_94_fu_3532_p2 = (z1_38_fu_3444_p3 ^ z0_37_fu_3338_p3);

assign xor_ln45_95_fu_3538_p2 = (z2_131_fu_3510_p3 ^ tmp_11_fu_3524_p3);

assign xor_ln45_98_fu_3604_p2 = (z1_35_fu_3252_p3 ^ z0_31_fu_2876_p3);

assign xor_ln45_99_fu_3610_p2 = (z2_132_fu_3556_p3 ^ tmp_13_fu_3596_p3);

assign xor_ln45_9_fu_582_p2 = (z2_121_fu_542_p3 ^ z0_1_fu_370_p3);

assign xor_ln45_fu_358_p2 = (z1_fu_346_p2 ^ z0_fu_328_p2);

assign z0_100_fu_9156_p2 = (b0_101_fu_9142_p2 & a0_309_fu_9128_p2);

assign z0_101_fu_9198_p3 = {{xor_ln45_256_fu_9186_p2}, {xor_ln45_257_fu_9192_p2}};

assign z0_102_fu_9262_p2 = (b0_102_fu_9248_p2 & a0_310_fu_9234_p2);

assign z0_103_fu_9328_p2 = (b0_103_fu_9220_p3 & a0_311_fu_9206_p3);

assign z0_104_fu_9460_p2 = (b0_105_fu_9072_p3 & a0_313_fu_9048_p3);

assign z0_105_fu_9502_p3 = {{xor_ln45_266_fu_9490_p2}, {xor_ln45_267_fu_9496_p2}};

assign z0_106_fu_9566_p2 = (b0_106_fu_9552_p2 & a0_314_fu_9538_p2);

assign z0_107_fu_9632_p2 = (b0_107_fu_9524_p3 & a0_315_fu_9510_p3);

assign z0_108_fu_9856_p2 = (b0_110_fu_8638_p3 & a0_318_fu_8588_p3);

assign z0_109_fu_9898_p3 = {{xor_ln45_280_fu_9886_p2}, {xor_ln45_281_fu_9892_p2}};

assign z0_10_fu_1050_p3 = {{xor_ln45_20_fu_1038_p2}, {xor_ln45_21_fu_1044_p2}};

assign z0_110_fu_9962_p2 = (b0_111_fu_9948_p2 & a0_319_fu_9934_p2);

assign z0_111_fu_10028_p2 = (b0_112_fu_9920_p3 & a0_320_fu_9906_p3);

assign z0_112_fu_10116_p3 = {{xor_ln45_288_fu_10104_p2}, {xor_ln45_289_fu_10110_p2}};

assign z0_113_fu_10232_p2 = (b0_114_fu_10218_p2 & a0_322_fu_10204_p2);

assign z0_114_fu_10274_p3 = {{xor_ln45_290_fu_10262_p2}, {xor_ln45_291_fu_10268_p2}};

assign z0_115_fu_10338_p2 = (b0_115_fu_10324_p2 & a0_323_fu_10310_p2);

assign z0_116_fu_10404_p2 = (b0_116_fu_10296_p3 & a0_324_fu_10282_p3);

assign z0_117_fu_10536_p2 = (b0_118_fu_10148_p3 & a0_326_fu_10124_p3);

assign z0_118_fu_10578_p3 = {{xor_ln45_300_fu_10566_p2}, {xor_ln45_301_fu_10572_p2}};

assign z0_119_fu_10642_p2 = (b0_119_fu_10628_p2 & a0_327_fu_10614_p2);

assign z0_11_fu_1114_p2 = (b0_13_fu_1100_p2 & a0_221_fu_1086_p2);

assign z0_120_fu_10708_p2 = (b0_120_fu_10600_p3 & a0_328_fu_10586_p3);

assign z0_12_fu_1180_p2 = (b0_14_fu_1072_p3 & a0_222_fu_1058_p3);

assign z0_13_fu_1340_p3 = {{xor_ln45_32_fu_1328_p2}, {xor_ln45_33_fu_1334_p2}};

assign z0_14_fu_1540_p2 = (b0_17_fu_1526_p2 & a0_225_fu_1512_p2);

assign z0_15_fu_1582_p3 = {{xor_ln45_34_fu_1570_p2}, {xor_ln45_35_fu_1576_p2}};

assign z0_16_fu_1646_p2 = (b0_18_fu_1632_p2 & a0_226_fu_1618_p2);

assign z0_17_fu_1712_p2 = (b0_19_fu_1604_p3 & a0_227_fu_1590_p3);

assign z0_18_fu_1800_p3 = {{xor_ln45_42_fu_1788_p2}, {xor_ln45_43_fu_1794_p2}};

assign z0_19_fu_1916_p2 = (b0_21_fu_1902_p2 & a0_229_fu_1888_p2);

assign z0_1_fu_370_p3 = {{xor_ln45_fu_358_p2}, {xor_ln45_1_fu_364_p2}};

assign z0_20_fu_1958_p3 = {{xor_ln45_44_fu_1946_p2}, {xor_ln45_45_fu_1952_p2}};

assign z0_21_fu_2022_p2 = (b0_22_fu_2008_p2 & a0_230_fu_1994_p2);

assign z0_22_fu_2088_p2 = (b0_23_fu_1980_p3 & a0_231_fu_1966_p3);

assign z0_23_fu_2220_p2 = (b0_25_fu_1832_p3 & a0_233_fu_1808_p3);

assign z0_24_fu_2262_p3 = {{xor_ln45_54_fu_2250_p2}, {xor_ln45_55_fu_2256_p2}};

assign z0_25_fu_2326_p2 = (b0_26_fu_2312_p2 & a0_234_fu_2298_p2);

assign z0_26_fu_2392_p2 = (b0_27_fu_2284_p3 & a0_235_fu_2270_p3);

assign z0_27_fu_2616_p2 = (b0_30_fu_1398_p3 & a0_238_fu_1348_p3);

assign z0_28_fu_2658_p3 = {{xor_ln45_68_fu_2646_p2}, {xor_ln45_69_fu_2652_p2}};

assign z0_29_fu_2722_p2 = (b0_31_fu_2708_p2 & a0_239_fu_2694_p2);

assign z0_2_fu_434_p2 = (b0_5_fu_420_p2 & a0_213_fu_406_p2);

assign z0_30_fu_2788_p2 = (b0_32_fu_2680_p3 & a0_240_fu_2666_p3);

assign z0_31_fu_2876_p3 = {{xor_ln45_76_fu_2864_p2}, {xor_ln45_77_fu_2870_p2}};

assign z0_32_fu_2992_p2 = (b0_34_fu_2978_p2 & a0_242_fu_2964_p2);

assign z0_33_fu_3034_p3 = {{xor_ln45_78_fu_3022_p2}, {xor_ln45_79_fu_3028_p2}};

assign z0_34_fu_3098_p2 = (b0_35_fu_3084_p2 & a0_243_fu_3070_p2);

assign z0_35_fu_3164_p2 = (b0_36_fu_3056_p3 & a0_244_fu_3042_p3);

assign z0_36_fu_3296_p2 = (b0_38_fu_2908_p3 & a0_246_fu_2884_p3);

assign z0_37_fu_3338_p3 = {{xor_ln45_88_fu_3326_p2}, {xor_ln45_89_fu_3332_p2}};

assign z0_38_fu_3402_p2 = (b0_39_fu_3388_p2 & a0_247_fu_3374_p2);

assign z0_39_fu_3468_p2 = (b0_40_fu_3360_p3 & a0_248_fu_3346_p3);

assign z0_3_fu_500_p2 = (b0_6_fu_392_p3 & a0_214_fu_378_p3);

assign z0_40_fu_3732_p3 = {{xor_ln45_104_fu_3720_p2}, {xor_ln45_105_fu_3726_p2}};

assign z0_41_fu_4080_p2 = (b0_44_fu_4066_p2 & a0_252_fu_4052_p2);

assign z0_42_fu_4122_p3 = {{xor_ln45_106_fu_4110_p2}, {xor_ln45_107_fu_4116_p2}};

assign z0_43_fu_4186_p2 = (b0_45_fu_4172_p2 & a0_253_fu_4158_p2);

assign z0_44_fu_4252_p2 = (b0_46_fu_4144_p3 & a0_254_fu_4130_p3);

assign z0_45_fu_4340_p3 = {{xor_ln45_114_fu_4328_p2}, {xor_ln45_115_fu_4334_p2}};

assign z0_46_fu_4456_p2 = (b0_48_fu_4442_p2 & a0_256_fu_4428_p2);

assign z0_47_fu_4498_p3 = {{xor_ln45_116_fu_4486_p2}, {xor_ln45_117_fu_4492_p2}};

assign z0_48_fu_4562_p2 = (b0_49_fu_4548_p2 & a0_257_fu_4534_p2);

assign z0_49_fu_4628_p2 = (b0_50_fu_4520_p3 & a0_258_fu_4506_p3);

assign z0_4_fu_588_p3 = {{xor_ln45_8_fu_576_p2}, {xor_ln45_9_fu_582_p2}};

assign z0_50_fu_4760_p2 = (b0_52_fu_4372_p3 & a0_260_fu_4348_p3);

assign z0_51_fu_4802_p3 = {{xor_ln45_126_fu_4790_p2}, {xor_ln45_127_fu_4796_p2}};

assign z0_52_fu_4866_p2 = (b0_53_fu_4852_p2 & a0_261_fu_4838_p2);

assign z0_53_fu_4932_p2 = (b0_54_fu_4824_p3 & a0_262_fu_4810_p3);

assign z0_54_fu_5092_p3 = {{xor_ln45_138_fu_5080_p2}, {xor_ln45_139_fu_5086_p2}};

assign z0_55_fu_5292_p2 = (b0_57_fu_5278_p2 & a0_265_fu_5264_p2);

assign z0_56_fu_5334_p3 = {{xor_ln45_140_fu_5322_p2}, {xor_ln45_141_fu_5328_p2}};

assign z0_57_fu_5398_p2 = (b0_58_fu_5384_p2 & a0_266_fu_5370_p2);

assign z0_58_fu_5464_p2 = (b0_59_fu_5356_p3 & a0_267_fu_5342_p3);

assign z0_59_fu_5552_p3 = {{xor_ln45_148_fu_5540_p2}, {xor_ln45_149_fu_5546_p2}};

assign z0_5_fu_704_p2 = (b0_8_fu_690_p2 & a0_216_fu_676_p2);

assign z0_60_fu_5668_p2 = (b0_61_fu_5654_p2 & a0_269_fu_5640_p2);

assign z0_61_fu_5710_p3 = {{xor_ln45_150_fu_5698_p2}, {xor_ln45_151_fu_5704_p2}};

assign z0_62_fu_5774_p2 = (b0_62_fu_5760_p2 & a0_270_fu_5746_p2);

assign z0_63_fu_5840_p2 = (b0_63_fu_5732_p3 & a0_271_fu_5718_p3);

assign z0_64_fu_5972_p2 = (b0_65_fu_5584_p3 & a0_273_fu_5560_p3);

assign z0_65_fu_6014_p3 = {{xor_ln45_160_fu_6002_p2}, {xor_ln45_161_fu_6008_p2}};

assign z0_66_fu_6078_p2 = (b0_66_fu_6064_p2 & a0_274_fu_6050_p2);

assign z0_67_fu_6144_p2 = (b0_67_fu_6036_p3 & a0_275_fu_6022_p3);

assign z0_68_fu_6368_p2 = (b0_70_fu_5150_p3 & a0_278_fu_5100_p3);

assign z0_69_fu_6410_p3 = {{xor_ln45_174_fu_6398_p2}, {xor_ln45_175_fu_6404_p2}};

assign z0_6_fu_746_p3 = {{xor_ln45_10_fu_734_p2}, {xor_ln45_11_fu_740_p2}};

assign z0_70_fu_6474_p2 = (b0_71_fu_6460_p2 & a0_279_fu_6446_p2);

assign z0_71_fu_6540_p2 = (b0_72_fu_6432_p3 & a0_280_fu_6418_p3);

assign z0_72_fu_6628_p3 = {{xor_ln45_182_fu_6616_p2}, {xor_ln45_183_fu_6622_p2}};

assign z0_73_fu_6744_p2 = (b0_74_fu_6730_p2 & a0_282_fu_6716_p2);

assign z0_74_fu_6786_p3 = {{xor_ln45_184_fu_6774_p2}, {xor_ln45_185_fu_6780_p2}};

assign z0_75_fu_6850_p2 = (b0_75_fu_6836_p2 & a0_283_fu_6822_p2);

assign z0_76_fu_6916_p2 = (b0_76_fu_6808_p3 & a0_284_fu_6794_p3);

assign z0_77_fu_7048_p2 = (b0_78_fu_6660_p3 & a0_286_fu_6636_p3);

assign z0_78_fu_7090_p3 = {{xor_ln45_194_fu_7078_p2}, {xor_ln45_195_fu_7084_p2}};

assign z0_79_fu_7154_p2 = (b0_79_fu_7140_p2 & a0_287_fu_7126_p2);

assign z0_7_fu_810_p2 = (b0_9_fu_796_p2 & a0_217_fu_782_p2);

assign z0_80_fu_7220_p2 = (b0_80_fu_7112_p3 & a0_288_fu_7098_p3);

assign z0_81_fu_7568_p2 = (b0_84_fu_3832_p3 & a0_292_fu_3740_p3);

assign z0_82_fu_7610_p3 = {{xor_ln45_212_fu_7598_p2}, {xor_ln45_213_fu_7604_p2}};

assign z0_83_fu_7674_p2 = (b0_85_fu_7660_p2 & a0_293_fu_7646_p2);

assign z0_84_fu_7740_p2 = (b0_86_fu_7632_p3 & a0_294_fu_7618_p3);

assign z0_85_fu_7828_p3 = {{xor_ln45_220_fu_7816_p2}, {xor_ln45_221_fu_7822_p2}};

assign z0_86_fu_7944_p2 = (b0_88_fu_7930_p2 & a0_296_fu_7916_p2);

assign z0_87_fu_7986_p3 = {{xor_ln45_222_fu_7974_p2}, {xor_ln45_223_fu_7980_p2}};

assign z0_88_fu_8050_p2 = (b0_89_fu_8036_p2 & a0_297_fu_8022_p2);

assign z0_89_fu_8116_p2 = (b0_90_fu_8008_p3 & a0_298_fu_7994_p3);

assign z0_8_fu_876_p2 = (b0_10_fu_768_p3 & a0_218_fu_754_p3);

assign z0_90_fu_8248_p2 = (b0_92_fu_7860_p3 & a0_300_fu_7836_p3);

assign z0_91_fu_8290_p3 = {{xor_ln45_232_fu_8278_p2}, {xor_ln45_233_fu_8284_p2}};

assign z0_92_fu_8354_p2 = (b0_93_fu_8340_p2 & a0_301_fu_8326_p2);

assign z0_93_fu_8420_p2 = (b0_94_fu_8312_p3 & a0_302_fu_8298_p3);

assign z0_94_fu_8580_p3 = {{xor_ln45_244_fu_8568_p2}, {xor_ln45_245_fu_8574_p2}};

assign z0_95_fu_8780_p2 = (b0_97_fu_8766_p2 & a0_305_fu_8752_p2);

assign z0_96_fu_8822_p3 = {{xor_ln45_246_fu_8810_p2}, {xor_ln45_247_fu_8816_p2}};

assign z0_97_fu_8886_p2 = (b0_98_fu_8872_p2 & a0_306_fu_8858_p2);

assign z0_98_fu_8952_p2 = (b0_99_fu_8844_p3 & a0_307_fu_8830_p3);

assign z0_99_fu_9040_p3 = {{xor_ln45_254_fu_9028_p2}, {xor_ln45_255_fu_9034_p2}};

assign z0_9_fu_1008_p2 = (b0_12_fu_620_p3 & a0_220_fu_596_p3);

assign z0_fu_328_p2 = (b0_4_fu_316_p1 & a0_212_fu_304_p1);

assign z1_100_fu_9304_p3 = {{xor_ln45_258_fu_9292_p2}, {xor_ln45_259_fu_9298_p2}};

assign z1_101_fu_9346_p2 = (b_309_fu_9340_p2 & a_351_fu_9334_p2);

assign z1_102_fu_9416_p3 = {{xor_ln45_264_fu_9404_p2}, {xor_ln45_265_fu_9410_p2}};

assign z1_103_fu_9478_p2 = (b_314_fu_9472_p2 & a_357_fu_9466_p2);

assign z1_104_fu_9584_p2 = (b_318_fu_9578_p2 & a_361_fu_9572_p2);

assign z1_105_fu_9608_p3 = {{xor_ln45_268_fu_9596_p2}, {xor_ln45_269_fu_9602_p2}};

assign z1_106_fu_9650_p2 = (b_322_fu_9644_p2 & a_365_fu_9638_p2);

assign z1_107_fu_9792_p3 = {{xor_ln45_278_fu_9780_p2}, {xor_ln45_279_fu_9786_p2}};

assign z1_108_fu_9874_p2 = (b_328_fu_9868_p2 & a_374_fu_9862_p2);

assign z1_109_fu_9980_p2 = (b_332_fu_9974_p2 & a_378_fu_9968_p2);

assign z1_10_fu_1132_p2 = (b_36_fu_1126_p2 & a_38_fu_1120_p2);

assign z1_110_fu_10004_p3 = {{xor_ln45_282_fu_9992_p2}, {xor_ln45_283_fu_9998_p2}};

assign z1_111_fu_10046_p2 = (b_336_fu_10040_p2 & a_382_fu_10034_p2);

assign z1_112_fu_10250_p2 = (b_341_fu_10244_p2 & a_388_fu_10238_p2);

assign z1_113_fu_10356_p2 = (b_345_fu_10350_p2 & a_392_fu_10344_p2);

assign z1_114_fu_10380_p3 = {{xor_ln45_292_fu_10368_p2}, {xor_ln45_293_fu_10374_p2}};

assign z1_115_fu_10422_p2 = (b_349_fu_10416_p2 & a_396_fu_10410_p2);

assign z1_116_fu_10492_p3 = {{xor_ln45_298_fu_10480_p2}, {xor_ln45_299_fu_10486_p2}};

assign z1_117_fu_10554_p2 = (b_354_fu_10548_p2 & a_402_fu_10542_p2);

assign z1_118_fu_10660_p2 = (b_358_fu_10654_p2 & a_406_fu_10648_p2);

assign z1_119_fu_10684_p3 = {{xor_ln45_302_fu_10672_p2}, {xor_ln45_303_fu_10678_p2}};

assign z1_11_fu_1156_p3 = {{xor_ln45_22_fu_1144_p2}, {xor_ln45_23_fu_1150_p2}};

assign z1_120_fu_10726_p2 = (b_362_fu_10720_p2 & a_410_fu_10714_p2);

assign z1_12_fu_1198_p2 = (b_40_fu_1192_p2 & a_42_fu_1186_p2);

assign z1_13_fu_1558_p2 = (b_46_fu_1552_p2 & a_51_fu_1546_p2);

assign z1_14_fu_1664_p2 = (b_50_fu_1658_p2 & a_55_fu_1652_p2);

assign z1_15_fu_1688_p3 = {{xor_ln45_36_fu_1676_p2}, {xor_ln45_37_fu_1682_p2}};

assign z1_16_fu_1730_p2 = (b_54_fu_1724_p2 & a_59_fu_1718_p2);

assign z1_17_fu_1934_p2 = (b_59_fu_1928_p2 & a_65_fu_1922_p2);

assign z1_18_fu_2040_p2 = (b_63_fu_2034_p2 & a_69_fu_2028_p2);

assign z1_19_fu_2064_p3 = {{xor_ln45_46_fu_2052_p2}, {xor_ln45_47_fu_2058_p2}};

assign z1_1_fu_452_p2 = (b_10_fu_446_p2 & a_10_fu_440_p2);

assign z1_20_fu_2106_p2 = (b_67_fu_2100_p2 & a_73_fu_2094_p2);

assign z1_21_fu_2176_p3 = {{xor_ln45_52_fu_2164_p2}, {xor_ln45_53_fu_2170_p2}};

assign z1_22_fu_2238_p2 = (b_72_fu_2232_p2 & a_79_fu_2226_p2);

assign z1_23_fu_2344_p2 = (b_76_fu_2338_p2 & a_83_fu_2332_p2);

assign z1_24_fu_2368_p3 = {{xor_ln45_56_fu_2356_p2}, {xor_ln45_57_fu_2362_p2}};

assign z1_25_fu_2410_p2 = (b_80_fu_2404_p2 & a_87_fu_2398_p2);

assign z1_26_fu_2552_p3 = {{xor_ln45_66_fu_2540_p2}, {xor_ln45_67_fu_2546_p2}};

assign z1_27_fu_2634_p2 = (b_86_fu_2628_p2 & a_96_fu_2622_p2);

assign z1_28_fu_2740_p2 = (b_90_fu_2734_p2 & a_100_fu_2728_p2);

assign z1_29_fu_2764_p3 = {{xor_ln45_70_fu_2752_p2}, {xor_ln45_71_fu_2758_p2}};

assign z1_2_fu_476_p3 = {{xor_ln45_2_fu_464_p2}, {xor_ln45_3_fu_470_p2}};

assign z1_30_fu_2806_p2 = (b_94_fu_2800_p2 & a_104_fu_2794_p2);

assign z1_31_fu_3010_p2 = (b_99_fu_3004_p2 & a_110_fu_2998_p2);

assign z1_32_fu_3116_p2 = (b_103_fu_3110_p2 & a_114_fu_3104_p2);

assign z1_33_fu_3140_p3 = {{xor_ln45_80_fu_3128_p2}, {xor_ln45_81_fu_3134_p2}};

assign z1_34_fu_3182_p2 = (b_107_fu_3176_p2 & a_118_fu_3170_p2);

assign z1_35_fu_3252_p3 = {{xor_ln45_86_fu_3240_p2}, {xor_ln45_87_fu_3246_p2}};

assign z1_36_fu_3314_p2 = (b_112_fu_3308_p2 & a_124_fu_3302_p2);

assign z1_37_fu_3420_p2 = (b_116_fu_3414_p2 & a_128_fu_3408_p2);

assign z1_38_fu_3444_p3 = {{xor_ln45_90_fu_3432_p2}, {xor_ln45_91_fu_3438_p2}};

assign z1_39_fu_3486_p2 = (b_120_fu_3480_p2 & a_132_fu_3474_p2);

assign z1_3_fu_518_p2 = (b_14_fu_512_p2 & a_14_fu_506_p2);

assign z1_40_fu_4098_p2 = (b_127_fu_4092_p2 & a_145_fu_4086_p2);

assign z1_41_fu_4204_p2 = (b_131_fu_4198_p2 & a_149_fu_4192_p2);

assign z1_42_fu_4228_p3 = {{xor_ln45_108_fu_4216_p2}, {xor_ln45_109_fu_4222_p2}};

assign z1_43_fu_4270_p2 = (b_135_fu_4264_p2 & a_153_fu_4258_p2);

assign z1_44_fu_4474_p2 = (b_140_fu_4468_p2 & a_159_fu_4462_p2);

assign z1_45_fu_4580_p2 = (b_144_fu_4574_p2 & a_163_fu_4568_p2);

assign z1_46_fu_4604_p3 = {{xor_ln45_118_fu_4592_p2}, {xor_ln45_119_fu_4598_p2}};

assign z1_47_fu_4646_p2 = (b_148_fu_4640_p2 & a_167_fu_4634_p2);

assign z1_48_fu_4716_p3 = {{xor_ln45_124_fu_4704_p2}, {xor_ln45_125_fu_4710_p2}};

assign z1_49_fu_4778_p2 = (b_153_fu_4772_p2 & a_173_fu_4766_p2);

assign z1_4_fu_722_p2 = (b_19_fu_716_p2 & a_20_fu_710_p2);

assign z1_50_fu_4884_p2 = (b_157_fu_4878_p2 & a_177_fu_4872_p2);

assign z1_51_fu_4908_p3 = {{xor_ln45_128_fu_4896_p2}, {xor_ln45_129_fu_4902_p2}};

assign z1_52_fu_4950_p2 = (b_161_fu_4944_p2 & a_181_fu_4938_p2);

assign z1_53_fu_5310_p2 = (b_167_fu_5304_p2 & a_190_fu_5298_p2);

assign z1_54_fu_5416_p2 = (b_171_fu_5410_p2 & a_194_fu_5404_p2);

assign z1_55_fu_5440_p3 = {{xor_ln45_142_fu_5428_p2}, {xor_ln45_143_fu_5434_p2}};

assign z1_56_fu_5482_p2 = (b_175_fu_5476_p2 & a_198_fu_5470_p2);

assign z1_57_fu_5686_p2 = (b_180_fu_5680_p2 & a_204_fu_5674_p2);

assign z1_58_fu_5792_p2 = (b_184_fu_5786_p2 & a_208_fu_5780_p2);

assign z1_59_fu_5816_p3 = {{xor_ln45_152_fu_5804_p2}, {xor_ln45_153_fu_5810_p2}};

assign z1_5_fu_828_p2 = (b_23_fu_822_p2 & a_24_fu_816_p2);

assign z1_60_fu_5858_p2 = (b_188_fu_5852_p2 & a_212_fu_5846_p2);

assign z1_61_fu_5928_p3 = {{xor_ln45_158_fu_5916_p2}, {xor_ln45_159_fu_5922_p2}};

assign z1_62_fu_5990_p2 = (b_193_fu_5984_p2 & a_218_fu_5978_p2);

assign z1_63_fu_6096_p2 = (b_197_fu_6090_p2 & a_222_fu_6084_p2);

assign z1_64_fu_6120_p3 = {{xor_ln45_162_fu_6108_p2}, {xor_ln45_163_fu_6114_p2}};

assign z1_65_fu_6162_p2 = (b_201_fu_6156_p2 & a_226_fu_6150_p2);

assign z1_66_fu_6304_p3 = {{xor_ln45_172_fu_6292_p2}, {xor_ln45_173_fu_6298_p2}};

assign z1_67_fu_6386_p2 = (b_207_fu_6380_p2 & a_235_fu_6374_p2);

assign z1_68_fu_6492_p2 = (b_211_fu_6486_p2 & a_239_fu_6480_p2);

assign z1_69_fu_6516_p3 = {{xor_ln45_176_fu_6504_p2}, {xor_ln45_177_fu_6510_p2}};

assign z1_6_fu_852_p3 = {{xor_ln45_12_fu_840_p2}, {xor_ln45_13_fu_846_p2}};

assign z1_70_fu_6558_p2 = (b_215_fu_6552_p2 & a_243_fu_6546_p2);

assign z1_71_fu_6762_p2 = (b_220_fu_6756_p2 & a_249_fu_6750_p2);

assign z1_72_fu_6868_p2 = (b_224_fu_6862_p2 & a_253_fu_6856_p2);

assign z1_73_fu_6892_p3 = {{xor_ln45_186_fu_6880_p2}, {xor_ln45_187_fu_6886_p2}};

assign z1_74_fu_6934_p2 = (b_228_fu_6928_p2 & a_257_fu_6922_p2);

assign z1_75_fu_7004_p3 = {{xor_ln45_192_fu_6992_p2}, {xor_ln45_193_fu_6998_p2}};

assign z1_76_fu_7066_p2 = (b_233_fu_7060_p2 & a_263_fu_7054_p2);

assign z1_77_fu_7172_p2 = (b_237_fu_7166_p2 & a_267_fu_7160_p2);

assign z1_78_fu_7196_p3 = {{xor_ln45_196_fu_7184_p2}, {xor_ln45_197_fu_7190_p2}};

assign z1_79_fu_7238_p2 = (b_241_fu_7232_p2 & a_271_fu_7226_p2);

assign z1_7_fu_894_p2 = (b_27_fu_888_p2 & a_28_fu_882_p2);

assign z1_80_fu_7484_p3 = {{xor_ln45_210_fu_7472_p2}, {xor_ln45_211_fu_7478_p2}};

assign z1_81_fu_7586_p2 = (b_248_fu_7580_p2 & a_284_fu_7574_p2);

assign z1_82_fu_7692_p2 = (b_252_fu_7686_p2 & a_288_fu_7680_p2);

assign z1_83_fu_7716_p3 = {{xor_ln45_214_fu_7704_p2}, {xor_ln45_215_fu_7710_p2}};

assign z1_84_fu_7758_p2 = (b_256_fu_7752_p2 & a_292_fu_7746_p2);

assign z1_85_fu_7962_p2 = (b_261_fu_7956_p2 & a_298_fu_7950_p2);

assign z1_86_fu_8068_p2 = (b_265_fu_8062_p2 & a_302_fu_8056_p2);

assign z1_87_fu_8092_p3 = {{xor_ln45_224_fu_8080_p2}, {xor_ln45_225_fu_8086_p2}};

assign z1_88_fu_8134_p2 = (b_269_fu_8128_p2 & a_306_fu_8122_p2);

assign z1_89_fu_8204_p3 = {{xor_ln45_230_fu_8192_p2}, {xor_ln45_231_fu_8198_p2}};

assign z1_8_fu_964_p3 = {{xor_ln45_18_fu_952_p2}, {xor_ln45_19_fu_958_p2}};

assign z1_90_fu_8266_p2 = (b_274_fu_8260_p2 & a_312_fu_8254_p2);

assign z1_91_fu_8372_p2 = (b_278_fu_8366_p2 & a_316_fu_8360_p2);

assign z1_92_fu_8396_p3 = {{xor_ln45_234_fu_8384_p2}, {xor_ln45_235_fu_8390_p2}};

assign z1_93_fu_8438_p2 = (b_282_fu_8432_p2 & a_320_fu_8426_p2);

assign z1_94_fu_8798_p2 = (b_288_fu_8792_p2 & a_329_fu_8786_p2);

assign z1_95_fu_8904_p2 = (b_292_fu_8898_p2 & a_333_fu_8892_p2);

assign z1_96_fu_8928_p3 = {{xor_ln45_248_fu_8916_p2}, {xor_ln45_249_fu_8922_p2}};

assign z1_97_fu_8970_p2 = (b_296_fu_8964_p2 & a_337_fu_8958_p2);

assign z1_98_fu_9174_p2 = (b_301_fu_9168_p2 & a_343_fu_9162_p2);

assign z1_99_fu_9280_p2 = (b_305_fu_9274_p2 & a_347_fu_9268_p2);

assign z1_9_fu_1026_p2 = (b_32_fu_1020_p2 & a_34_fu_1014_p2);

assign z1_fu_346_p2 = (b_6_fu_340_p2 & a_6_fu_334_p2);

assign z2_101_fu_9484_p2 = (b1_221_fu_9452_p3 & a1_321_fu_9444_p3);

assign z2_102_fu_9590_p2 = (b1_222_fu_9558_p3 & a1_322_fu_9544_p3);

assign z2_103_fu_9656_p2 = (b1_223_fu_9624_p3 & a1_323_fu_9616_p3);

assign z2_106_fu_9880_p2 = (b1_226_fu_9848_p3 & a1_327_fu_9840_p3);

assign z2_107_fu_9986_p2 = (b1_227_fu_9954_p3 & a1_328_fu_9940_p3);

assign z2_108_fu_10052_p2 = (b1_228_fu_10020_p3 & a1_329_fu_10012_p3);

assign z2_10_fu_1204_p2 = (b1_130_fu_1172_p3 & a1_219_fu_1164_p3);

assign z2_110_fu_10256_p2 = (b1_230_fu_10224_p3 & a1_331_fu_10210_p3);

assign z2_111_fu_10362_p2 = (b1_231_fu_10330_p3 & a1_332_fu_10316_p3);

assign z2_112_fu_10428_p2 = (b1_232_fu_10396_p3 & a1_333_fu_10388_p3);

assign z2_114_fu_10560_p2 = (b1_234_fu_10528_p3 & a1_335_fu_10520_p3);

assign z2_115_fu_10666_p2 = (b1_235_fu_10634_p3 & a1_336_fu_10620_p3);

assign z2_116_fu_10732_p2 = (b1_236_fu_10700_p3 & a1_337_fu_10692_p3);

assign z2_121_fu_542_p3 = {{a1_9_fu_530_p2}, {a0_fu_536_p2}};

assign z2_122_fu_918_p3 = {{a1_15_fu_906_p2}, {a0_13_fu_912_p2}};

assign z2_123_fu_1222_p3 = {{a1_21_fu_1210_p2}, {a0_20_fu_1216_p2}};

assign z2_124_fu_1268_p3 = {{a1_220_fu_1256_p2}, {a0_21_fu_1262_p2}};

assign z2_125_fu_1754_p3 = {{a1_31_fu_1742_p2}, {a0_32_fu_1748_p2}};

assign z2_126_fu_2130_p3 = {{a1_37_fu_2118_p2}, {a0_39_fu_2124_p2}};

assign z2_127_fu_2434_p3 = {{a1_42_fu_2422_p2}, {a0_46_fu_2428_p2}};

assign z2_128_fu_2480_p3 = {{a1_234_fu_2468_p2}, {a0_47_fu_2474_p2}};

assign z2_129_fu_2830_p3 = {{a1_52_fu_2818_p2}, {a0_54_fu_2824_p2}};

assign z2_130_fu_3206_p3 = {{a1_58_fu_3194_p2}, {a0_62_fu_3200_p2}};

assign z2_131_fu_3510_p3 = {{a1_63_fu_3498_p2}, {a0_69_fu_3504_p2}};

assign z2_132_fu_3556_p3 = {{a1_248_fu_3544_p2}, {a0_72_fu_3550_p2}};

assign z2_133_fu_3628_p3 = {{a1_249_fu_3616_p2}, {a0_75_fu_3622_p2}};

assign z2_134_fu_4294_p3 = {{a1_78_fu_4282_p2}, {a0_90_fu_4288_p2}};

assign z2_135_fu_4670_p3 = {{a1_84_fu_4658_p2}, {a0_97_fu_4664_p2}};

assign z2_136_fu_4974_p3 = {{a1_90_fu_4962_p2}, {a0_102_fu_4968_p2}};

assign z2_137_fu_5020_p3 = {{a1_265_fu_5008_p2}, {a0_103_fu_5014_p2}};

assign z2_138_fu_5506_p3 = {{a1_99_fu_5494_p2}, {a0_114_fu_5500_p2}};

assign z2_139_fu_5882_p3 = {{a1_105_fu_5870_p2}, {a0_123_fu_5876_p2}};

assign z2_13_fu_1564_p2 = (b1_133_fu_1532_p3 & a1_223_fu_1518_p3);

assign z2_140_fu_6186_p3 = {{a1_112_fu_6174_p2}, {a0_129_fu_6180_p2}};

assign z2_141_fu_6232_p3 = {{a1_279_fu_6220_p2}, {a0_130_fu_6226_p2}};

assign z2_142_fu_6582_p3 = {{a1_120_fu_6570_p2}, {a0_135_fu_6576_p2}};

assign z2_143_fu_6958_p3 = {{a1_126_fu_6946_p2}, {a0_140_fu_6952_p2}};

assign z2_144_fu_7262_p3 = {{a1_133_fu_7250_p2}, {a0_144_fu_7256_p2}};

assign z2_145_fu_7308_p3 = {{a1_293_fu_7296_p2}, {a0_145_fu_7302_p2}};

assign z2_146_fu_7380_p3 = {{a1_294_fu_7368_p2}, {a0_147_fu_7374_p2}};

assign z2_147_fu_7782_p3 = {{a1_147_fu_7770_p2}, {a0_154_fu_7776_p2}};

assign z2_148_fu_8158_p3 = {{a1_153_fu_8146_p2}, {a0_159_fu_8152_p2}};

assign z2_149_fu_8462_p3 = {{a1_159_fu_8450_p2}, {a0_164_fu_8456_p2}};

assign z2_14_fu_1670_p2 = (b1_134_fu_1638_p3 & a1_224_fu_1624_p3);

assign z2_150_fu_8508_p3 = {{a1_310_fu_8496_p2}, {a0_165_fu_8502_p2}};

assign z2_151_fu_8994_p3 = {{a1_168_fu_8982_p2}, {a0_172_fu_8988_p2}};

assign z2_152_fu_9370_p3 = {{a1_173_fu_9358_p2}, {a0_177_fu_9364_p2}};

assign z2_153_fu_9674_p3 = {{a1_178_fu_9662_p2}, {a0_181_fu_9668_p2}};

assign z2_154_fu_9720_p3 = {{a1_324_fu_9708_p2}, {a0_182_fu_9714_p2}};

assign z2_155_fu_10070_p3 = {{a1_186_fu_10058_p2}, {a0_188_fu_10064_p2}};

assign z2_156_fu_10446_p3 = {{a1_191_fu_10434_p2}, {a0_193_fu_10440_p2}};

assign z2_157_fu_10750_p3 = {{a1_fu_10738_p2}, {a0_198_fu_10744_p2}};

assign z2_158_fu_10796_p3 = {{a1_338_fu_10784_p2}, {a0_199_fu_10790_p2}};

assign z2_159_fu_10868_p3 = {{a1_339_fu_10856_p2}, {a0_201_fu_10862_p2}};

assign z2_15_fu_1736_p2 = (b1_135_fu_1704_p3 & a1_225_fu_1696_p3);

assign z2_160_fu_10972_p3 = {{a1_341_fu_10960_p2}, {a0_204_fu_10966_p2}};

assign z2_17_fu_1940_p2 = (b1_137_fu_1908_p3 & a1_227_fu_1894_p3);

assign z2_18_fu_2046_p2 = (b1_138_fu_2014_p3 & a1_228_fu_2000_p3);

assign z2_19_fu_2112_p2 = (b1_139_fu_2080_p3 & a1_229_fu_2072_p3);

assign z2_1_fu_458_p2 = (b1_121_fu_426_p3 & a1_210_fu_412_p3);

assign z2_21_fu_2244_p2 = (b1_141_fu_2212_p3 & a1_231_fu_2204_p3);

assign z2_22_fu_2350_p2 = (b1_142_fu_2318_p3 & a1_232_fu_2304_p3);

assign z2_23_fu_2416_p2 = (b1_143_fu_2384_p3 & a1_233_fu_2376_p3);

assign z2_26_fu_2640_p2 = (b1_146_fu_2608_p3 & a1_237_fu_2600_p3);

assign z2_27_fu_2746_p2 = (b1_147_fu_2714_p3 & a1_238_fu_2700_p3);

assign z2_28_fu_2812_p2 = (b1_148_fu_2780_p3 & a1_239_fu_2772_p3);

assign z2_2_fu_524_p2 = (b1_122_fu_492_p3 & a1_211_fu_484_p3);

assign z2_30_fu_3016_p2 = (b1_150_fu_2984_p3 & a1_241_fu_2970_p3);

assign z2_31_fu_3122_p2 = (b1_151_fu_3090_p3 & a1_242_fu_3076_p3);

assign z2_32_fu_3188_p2 = (b1_152_fu_3156_p3 & a1_243_fu_3148_p3);

assign z2_34_fu_3320_p2 = (b1_154_fu_3288_p3 & a1_245_fu_3280_p3);

assign z2_35_fu_3426_p2 = (b1_155_fu_3394_p3 & a1_246_fu_3380_p3);

assign z2_36_fu_3492_p2 = (b1_156_fu_3460_p3 & a1_247_fu_3452_p3);

assign z2_40_fu_4104_p2 = (b1_160_fu_4072_p3 & a1_254_fu_4058_p3);

assign z2_41_fu_4210_p2 = (b1_161_fu_4178_p3 & a1_255_fu_4164_p3);

assign z2_42_fu_4276_p2 = (b1_162_fu_4244_p3 & a1_256_fu_4236_p3);

assign z2_44_fu_4480_p2 = (b1_164_fu_4448_p3 & a1_258_fu_4434_p3);

assign z2_45_fu_4586_p2 = (b1_165_fu_4554_p3 & a1_259_fu_4540_p3);

assign z2_46_fu_4652_p2 = (b1_166_fu_4620_p3 & a1_260_fu_4612_p3);

assign z2_48_fu_4784_p2 = (b1_168_fu_4752_p3 & a1_262_fu_4744_p3);

assign z2_49_fu_4890_p2 = (b1_169_fu_4858_p3 & a1_263_fu_4844_p3);

assign z2_4_fu_728_p2 = (b1_124_fu_696_p3 & a1_213_fu_682_p3);

assign z2_50_fu_4956_p2 = (b1_170_fu_4924_p3 & a1_264_fu_4916_p3);

assign z2_53_fu_5316_p2 = (b1_173_fu_5284_p3 & a1_268_fu_5270_p3);

assign z2_54_fu_5422_p2 = (b1_174_fu_5390_p3 & a1_269_fu_5376_p3);

assign z2_55_fu_5488_p2 = (b1_175_fu_5456_p3 & a1_270_fu_5448_p3);

assign z2_57_fu_5692_p2 = (b1_177_fu_5660_p3 & a1_272_fu_5646_p3);

assign z2_58_fu_5798_p2 = (b1_178_fu_5766_p3 & a1_273_fu_5752_p3);

assign z2_59_fu_5864_p2 = (b1_179_fu_5832_p3 & a1_274_fu_5824_p3);

assign z2_5_fu_834_p2 = (b1_125_fu_802_p3 & a1_214_fu_788_p3);

assign z2_61_fu_5996_p2 = (b1_181_fu_5964_p3 & a1_276_fu_5956_p3);

assign z2_62_fu_6102_p2 = (b1_182_fu_6070_p3 & a1_277_fu_6056_p3);

assign z2_63_fu_6168_p2 = (b1_183_fu_6136_p3 & a1_278_fu_6128_p3);

assign z2_66_fu_6392_p2 = (b1_186_fu_6360_p3 & a1_282_fu_6352_p3);

assign z2_67_fu_6498_p2 = (b1_187_fu_6466_p3 & a1_283_fu_6452_p3);

assign z2_68_fu_6564_p2 = (b1_188_fu_6532_p3 & a1_284_fu_6524_p3);

assign z2_6_fu_900_p2 = (b1_126_fu_868_p3 & a1_215_fu_860_p3);

assign z2_70_fu_6768_p2 = (b1_190_fu_6736_p3 & a1_286_fu_6722_p3);

assign z2_71_fu_6874_p2 = (b1_191_fu_6842_p3 & a1_287_fu_6828_p3);

assign z2_72_fu_6940_p2 = (b1_192_fu_6908_p3 & a1_288_fu_6900_p3);

assign z2_74_fu_7072_p2 = (b1_194_fu_7040_p3 & a1_290_fu_7032_p3);

assign z2_75_fu_7178_p2 = (b1_195_fu_7146_p3 & a1_291_fu_7132_p3);

assign z2_76_fu_7244_p2 = (b1_196_fu_7212_p3 & a1_292_fu_7204_p3);

assign z2_80_fu_7592_p2 = (b1_200_fu_7560_p3 & a1_299_fu_7552_p3);

assign z2_81_fu_7698_p2 = (b1_201_fu_7666_p3 & a1_300_fu_7652_p3);

assign z2_82_fu_7764_p2 = (b1_202_fu_7732_p3 & a1_301_fu_7724_p3);

assign z2_84_fu_7968_p2 = (b1_204_fu_7936_p3 & a1_303_fu_7922_p3);

assign z2_85_fu_8074_p2 = (b1_205_fu_8042_p3 & a1_304_fu_8028_p3);

assign z2_86_fu_8140_p2 = (b1_206_fu_8108_p3 & a1_305_fu_8100_p3);

assign z2_88_fu_8272_p2 = (b1_208_fu_8240_p3 & a1_307_fu_8232_p3);

assign z2_89_fu_8378_p2 = (b1_209_fu_8346_p3 & a1_308_fu_8332_p3);

assign z2_8_fu_1032_p2 = (b1_128_fu_1000_p3 & a1_217_fu_992_p3);

assign z2_90_fu_8444_p2 = (b1_210_fu_8412_p3 & a1_309_fu_8404_p3);

assign z2_93_fu_8804_p2 = (b1_213_fu_8772_p3 & a1_313_fu_8758_p3);

assign z2_94_fu_8910_p2 = (b1_214_fu_8878_p3 & a1_314_fu_8864_p3);

assign z2_95_fu_8976_p2 = (b1_215_fu_8944_p3 & a1_315_fu_8936_p3);

assign z2_97_fu_9180_p2 = (b1_217_fu_9148_p3 & a1_317_fu_9134_p3);

assign z2_98_fu_9286_p2 = (b1_218_fu_9254_p3 & a1_318_fu_9240_p3);

assign z2_99_fu_9352_p2 = (b1_219_fu_9320_p3 & a1_319_fu_9312_p3);

assign z2_9_fu_1138_p2 = (b1_129_fu_1106_p3 & a1_218_fu_1092_p3);

assign z2_fu_352_p2 = (b1_120_fu_320_p3 & a1_209_fu_308_p3);

assign ap_return = {{xor_ln45_320_fu_11098_p2}, {xor_ln45_321_fu_11104_p2}};

endmodule //binary_tower_32b_mul
