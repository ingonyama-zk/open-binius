module binary_tower_32b_mul (
        input ap_clk,
        input ap_rst,
        input ap_ce,
        input  [31:0] a,
        input  [31:0] b,
        output [31:0] ap_return
);

wire   [0:0] trunc_ln86_fu_214_p1;
wire   [0:0] trunc_ln86_1_fu_218_p1;
wire   [0:0] tmp_fu_228_p3;
wire   [0:0] tmp_1_fu_236_p3;
wire   [0:0] tmp_2_fu_250_p3;
wire   [0:0] tmp_3_fu_258_p3;
wire   [0:0] tmp_4_fu_272_p3;
wire   [0:0] tmp_5_fu_280_p3;
wire   [0:0] and_ln86_fu_222_p2;
wire   [0:0] and_ln86_1_fu_244_p2;
wire   [0:0] and_ln86_2_fu_266_p2;
wire   [0:0] and_ln86_3_fu_288_p2;
wire   [0:0] xor_ln86_1_fu_300_p2;
wire   [0:0] xor_ln86_fu_294_p2;
wire   [0:0] and_ln87_1_fu_318_p2;
wire   [0:0] xor_ln87_fu_336_p2;
wire   [0:0] and_ln87_fu_312_p2;
wire   [0:0] and_ln87_3_fu_330_p2;
wire   [0:0] xor_ln87_2_fu_348_p2;
wire   [0:0] and_ln87_2_fu_324_p2;
wire   [0:0] xor_ln87_3_fu_354_p2;
wire   [0:0] xor_ln87_1_fu_342_p2;
wire   [0:0] and_ln88_1_fu_372_p2;
wire   [0:0] and_ln88_2_fu_378_p2;
wire   [0:0] xor_ln88_fu_390_p2;
wire   [0:0] and_ln88_fu_366_p2;
wire   [0:0] and_ln88_3_fu_384_p2;
wire   [0:0] xor_ln88_2_fu_402_p2;
wire   [0:0] xor_ln88_3_fu_408_p2;
wire   [0:0] xor_ln88_1_fu_396_p2;
wire   [0:0] and_ln90_fu_420_p2;
wire   [0:0] and_ln90_1_fu_426_p2;
wire   [0:0] and_ln90_2_fu_432_p2;
wire   [0:0] xor_ln91_2_fu_450_p2;
wire   [0:0] xor_ln91_fu_444_p2;
wire   [0:0] xor_ln91_8_fu_468_p2;
wire   [0:0] and_ln91_fu_438_p2;
wire   [0:0] xor_ln91_10_fu_474_p2;
wire   [0:0] xor_ln91_6_fu_462_p2;
wire   [0:0] xor_ln91_12_fu_480_p2;
wire   [0:0] xor_ln91_4_fu_456_p2;
wire   [0:0] xor_ln91_1_fu_486_p2;
wire   [0:0] xor_ln88_4_fu_414_p2;
wire   [0:0] xor_ln87_4_fu_360_p2;
wire   [0:0] xor_ln86_2_fu_306_p2;
wire   [3:0] a1_12_fu_190_p4;
wire   [3:0] a0_13_fu_186_p1;
wire   [3:0] b1_12_fu_204_p4;
wire   [3:0] b0_2_fu_200_p1;
wire   [3:0] a_4_fu_504_p2;
wire   [3:0] b_4_fu_510_p2;
wire   [0:0] trunc_ln86_2_fu_516_p1;
wire   [0:0] trunc_ln86_3_fu_520_p1;
wire   [0:0] tmp_6_fu_530_p3;
wire   [0:0] tmp_7_fu_538_p3;
wire   [0:0] tmp_8_fu_552_p3;
wire   [0:0] tmp_9_fu_560_p3;
wire   [0:0] tmp_10_fu_574_p3;
wire   [0:0] tmp_11_fu_582_p3;
wire   [0:0] and_ln86_4_fu_524_p2;
wire   [0:0] and_ln86_5_fu_546_p2;
wire   [0:0] and_ln86_6_fu_568_p2;
wire   [0:0] and_ln86_7_fu_590_p2;
wire   [0:0] xor_ln86_4_fu_602_p2;
wire   [0:0] xor_ln86_3_fu_596_p2;
wire   [0:0] and_ln87_5_fu_620_p2;
wire   [0:0] xor_ln87_5_fu_638_p2;
wire   [0:0] and_ln87_4_fu_614_p2;
wire   [0:0] and_ln87_7_fu_632_p2;
wire   [0:0] xor_ln87_7_fu_650_p2;
wire   [0:0] and_ln87_6_fu_626_p2;
wire   [0:0] xor_ln87_8_fu_656_p2;
wire   [0:0] xor_ln87_6_fu_644_p2;
wire   [0:0] and_ln88_5_fu_674_p2;
wire   [0:0] and_ln88_6_fu_680_p2;
wire   [0:0] xor_ln88_5_fu_692_p2;
wire   [0:0] and_ln88_4_fu_668_p2;
wire   [0:0] and_ln88_7_fu_686_p2;
wire   [0:0] xor_ln88_7_fu_704_p2;
wire   [0:0] xor_ln88_8_fu_710_p2;
wire   [0:0] xor_ln88_6_fu_698_p2;
wire   [0:0] and_ln90_3_fu_722_p2;
wire   [0:0] and_ln90_4_fu_728_p2;
wire   [0:0] and_ln90_5_fu_734_p2;
wire   [0:0] xor_ln91_16_fu_752_p2;
wire   [0:0] xor_ln91_14_fu_746_p2;
wire   [0:0] xor_ln91_22_fu_770_p2;
wire   [0:0] and_ln91_1_fu_740_p2;
wire   [0:0] xor_ln91_24_fu_776_p2;
wire   [0:0] xor_ln91_20_fu_764_p2;
wire   [0:0] xor_ln91_26_fu_782_p2;
wire   [0:0] xor_ln91_18_fu_758_p2;
wire   [0:0] xor_ln91_3_fu_788_p2;
wire   [0:0] xor_ln88_9_fu_716_p2;
wire   [0:0] xor_ln87_9_fu_662_p2;
wire   [0:0] xor_ln86_5_fu_608_p2;
wire   [0:0] tmp_12_fu_806_p3;
wire   [0:0] tmp_13_fu_814_p3;
wire   [0:0] tmp_14_fu_828_p3;
wire   [0:0] tmp_15_fu_836_p3;
wire   [0:0] tmp_16_fu_850_p3;
wire   [0:0] tmp_17_fu_858_p3;
wire   [0:0] tmp_18_fu_872_p3;
wire   [0:0] tmp_19_fu_880_p3;
wire   [0:0] and_ln86_9_fu_844_p2;
wire   [0:0] and_ln86_10_fu_866_p2;
wire   [0:0] and_ln86_8_fu_822_p2;
wire   [0:0] and_ln86_11_fu_888_p2;
wire   [0:0] xor_ln86_7_fu_900_p2;
wire   [0:0] xor_ln86_6_fu_894_p2;
wire   [0:0] and_ln87_9_fu_918_p2;
wire   [0:0] and_ln87_8_fu_912_p2;
wire   [0:0] and_ln87_10_fu_924_p2;
wire   [0:0] xor_ln87_11_fu_936_p2;
wire   [0:0] xor_ln87_10_fu_930_p2;
wire   [0:0] and_ln87_11_fu_948_p2;
wire   [0:0] xor_ln87_13_fu_954_p2;
wire   [0:0] xor_ln87_12_fu_942_p2;
wire   [0:0] and_ln88_10_fu_978_p2;
wire   [0:0] and_ln88_8_fu_966_p2;
wire   [0:0] and_ln88_11_fu_984_p2;
wire   [0:0] xor_ln88_11_fu_996_p2;
wire   [0:0] and_ln88_9_fu_972_p2;
wire   [0:0] xor_ln88_12_fu_1002_p2;
wire   [0:0] xor_ln88_10_fu_990_p2;
wire   [0:0] xor_ln88_13_fu_1008_p2;
wire   [0:0] and_ln91_2_fu_1038_p2;
wire   [0:0] xor_ln91_30_fu_1050_p2;
wire   [0:0] xor_ln91_28_fu_1044_p2;
wire   [0:0] and_ln90_7_fu_1026_p2;
wire   [0:0] and_ln90_6_fu_1020_p2;
wire   [0:0] xor_ln91_36_fu_1068_p2;
wire   [0:0] and_ln90_8_fu_1032_p2;
wire   [0:0] xor_ln91_38_fu_1074_p2;
wire   [0:0] xor_ln91_34_fu_1062_p2;
wire   [0:0] xor_ln91_40_fu_1080_p2;
wire   [0:0] xor_ln91_32_fu_1056_p2;
wire   [0:0] xor_ln91_5_fu_1086_p2;
wire   [0:0] xor_ln88_14_fu_1014_p2;
wire   [0:0] xor_ln87_14_fu_960_p2;
wire   [0:0] xor_ln86_8_fu_906_p2;
wire   [0:0] xor_ln54_fu_1110_p2;
wire   [0:0] xor_ln54_1_fu_1116_p2;
wire   [0:0] xor_ln53_fu_1104_p2;
wire   [3:0] res_41_fu_794_p5;
wire   [3:0] res_40_fu_492_p5;
wire   [3:0] res_42_fu_1092_p5;
wire   [3:0] res_fu_1122_p5;
wire   [3:0] xor_ln101_1_fu_1140_p2;
wire   [3:0] xor_ln101_fu_1134_p2;
wire   [3:0] xor_ln101_2_fu_1146_p2;
wire   [3:0] xor_ln101_3_fu_1152_p2;
wire   [7:0] a1_11_fu_162_p4;
wire   [7:0] a0_12_fu_158_p1;
wire   [7:0] b1_11_fu_176_p4;
wire   [7:0] b0_1_fu_172_p1;
wire   [7:0] a_7_fu_1176_p2;
wire   [7:0] b_6_fu_1192_p2;
wire   [0:0] trunc_ln86_4_fu_1218_p1;
wire   [0:0] trunc_ln86_5_fu_1222_p1;
wire   [0:0] tmp_20_fu_1232_p3;
wire   [0:0] tmp_21_fu_1240_p3;
wire   [0:0] tmp_22_fu_1254_p3;
wire   [0:0] tmp_23_fu_1262_p3;
wire   [0:0] tmp_24_fu_1276_p3;
wire   [0:0] tmp_25_fu_1284_p3;
wire   [0:0] and_ln86_12_fu_1226_p2;
wire   [0:0] and_ln86_13_fu_1248_p2;
wire   [0:0] and_ln86_14_fu_1270_p2;
wire   [0:0] and_ln86_15_fu_1292_p2;
wire   [0:0] xor_ln86_10_fu_1304_p2;
wire   [0:0] xor_ln86_9_fu_1298_p2;
wire   [0:0] and_ln87_13_fu_1322_p2;
wire   [0:0] xor_ln87_15_fu_1340_p2;
wire   [0:0] and_ln87_12_fu_1316_p2;
wire   [0:0] and_ln87_15_fu_1334_p2;
wire   [0:0] xor_ln87_17_fu_1352_p2;
wire   [0:0] and_ln87_14_fu_1328_p2;
wire   [0:0] xor_ln87_18_fu_1358_p2;
wire   [0:0] xor_ln87_16_fu_1346_p2;
wire   [0:0] and_ln88_13_fu_1376_p2;
wire   [0:0] and_ln88_14_fu_1382_p2;
wire   [0:0] xor_ln88_15_fu_1394_p2;
wire   [0:0] and_ln88_12_fu_1370_p2;
wire   [0:0] and_ln88_15_fu_1388_p2;
wire   [0:0] xor_ln88_17_fu_1406_p2;
wire   [0:0] xor_ln88_18_fu_1412_p2;
wire   [0:0] xor_ln88_16_fu_1400_p2;
wire   [0:0] and_ln90_9_fu_1424_p2;
wire   [0:0] and_ln90_10_fu_1430_p2;
wire   [0:0] and_ln90_11_fu_1436_p2;
wire   [0:0] xor_ln91_44_fu_1454_p2;
wire   [0:0] xor_ln91_42_fu_1448_p2;
wire   [0:0] xor_ln91_50_fu_1472_p2;
wire   [0:0] and_ln91_3_fu_1442_p2;
wire   [0:0] xor_ln91_52_fu_1478_p2;
wire   [0:0] xor_ln91_48_fu_1466_p2;
wire   [0:0] xor_ln91_54_fu_1484_p2;
wire   [0:0] xor_ln91_46_fu_1460_p2;
wire   [0:0] xor_ln91_7_fu_1490_p2;
wire   [0:0] xor_ln88_19_fu_1418_p2;
wire   [0:0] xor_ln87_19_fu_1364_p2;
wire   [0:0] xor_ln86_11_fu_1310_p2;
wire   [3:0] a1_13_fu_1198_p4;
wire   [3:0] xor_ln99_fu_1508_p2;
wire   [3:0] a0_14_fu_1166_p4;
wire   [3:0] b1_13_fu_1208_p4;
wire   [3:0] xor_ln99_4_fu_1520_p2;
wire   [3:0] b0_3_fu_1182_p4;
wire   [3:0] a_8_fu_1514_p2;
wire   [3:0] b_7_fu_1526_p2;
wire   [0:0] trunc_ln86_6_fu_1532_p1;
wire   [0:0] trunc_ln86_7_fu_1536_p1;
wire   [0:0] tmp_26_fu_1546_p3;
wire   [0:0] tmp_27_fu_1554_p3;
wire   [0:0] tmp_28_fu_1568_p3;
wire   [0:0] tmp_29_fu_1576_p3;
wire   [0:0] tmp_30_fu_1590_p3;
wire   [0:0] tmp_31_fu_1598_p3;
wire   [0:0] and_ln86_16_fu_1540_p2;
wire   [0:0] and_ln86_17_fu_1562_p2;
wire   [0:0] and_ln86_18_fu_1584_p2;
wire   [0:0] and_ln86_19_fu_1606_p2;
wire   [0:0] xor_ln86_13_fu_1618_p2;
wire   [0:0] xor_ln86_12_fu_1612_p2;
wire   [0:0] and_ln87_17_fu_1636_p2;
wire   [0:0] xor_ln87_20_fu_1654_p2;
wire   [0:0] and_ln87_16_fu_1630_p2;
wire   [0:0] and_ln87_19_fu_1648_p2;
wire   [0:0] xor_ln87_22_fu_1666_p2;
wire   [0:0] and_ln87_18_fu_1642_p2;
wire   [0:0] xor_ln87_23_fu_1672_p2;
wire   [0:0] xor_ln87_21_fu_1660_p2;
wire   [0:0] and_ln88_17_fu_1690_p2;
wire   [0:0] and_ln88_18_fu_1696_p2;
wire   [0:0] xor_ln88_20_fu_1708_p2;
wire   [0:0] and_ln88_16_fu_1684_p2;
wire   [0:0] and_ln88_19_fu_1702_p2;
wire   [0:0] xor_ln88_22_fu_1720_p2;
wire   [0:0] xor_ln88_23_fu_1726_p2;
wire   [0:0] xor_ln88_21_fu_1714_p2;
wire   [0:0] and_ln90_12_fu_1738_p2;
wire   [0:0] and_ln90_13_fu_1744_p2;
wire   [0:0] and_ln90_14_fu_1750_p2;
wire   [0:0] xor_ln91_56_fu_1768_p2;
wire   [0:0] xor_ln91_55_fu_1762_p2;
wire   [0:0] xor_ln91_59_fu_1786_p2;
wire   [0:0] and_ln91_4_fu_1756_p2;
wire   [0:0] xor_ln91_60_fu_1792_p2;
wire   [0:0] xor_ln91_58_fu_1780_p2;
wire   [0:0] xor_ln91_61_fu_1798_p2;
wire   [0:0] xor_ln91_57_fu_1774_p2;
wire   [0:0] xor_ln91_9_fu_1804_p2;
wire   [0:0] xor_ln88_24_fu_1732_p2;
wire   [0:0] xor_ln87_24_fu_1678_p2;
wire   [0:0] xor_ln86_14_fu_1624_p2;
wire   [0:0] tmp_32_fu_1822_p3;
wire   [0:0] tmp_33_fu_1830_p3;
wire   [0:0] tmp_34_fu_1844_p3;
wire   [0:0] tmp_35_fu_1852_p3;
wire   [0:0] tmp_36_fu_1866_p3;
wire   [0:0] tmp_37_fu_1874_p3;
wire   [0:0] tmp_38_fu_1888_p3;
wire   [0:0] tmp_39_fu_1896_p3;
wire   [0:0] and_ln86_21_fu_1860_p2;
wire   [0:0] and_ln86_22_fu_1882_p2;
wire   [0:0] and_ln86_20_fu_1838_p2;
wire   [0:0] and_ln86_23_fu_1904_p2;
wire   [0:0] xor_ln86_16_fu_1916_p2;
wire   [0:0] xor_ln86_15_fu_1910_p2;
wire   [0:0] and_ln87_21_fu_1934_p2;
wire   [0:0] and_ln87_20_fu_1928_p2;
wire   [0:0] and_ln87_22_fu_1940_p2;
wire   [0:0] xor_ln87_26_fu_1952_p2;
wire   [0:0] xor_ln87_25_fu_1946_p2;
wire   [0:0] and_ln87_23_fu_1964_p2;
wire   [0:0] xor_ln87_28_fu_1970_p2;
wire   [0:0] xor_ln87_27_fu_1958_p2;
wire   [0:0] and_ln88_22_fu_1994_p2;
wire   [0:0] and_ln88_20_fu_1982_p2;
wire   [0:0] and_ln88_23_fu_2000_p2;
wire   [0:0] xor_ln88_26_fu_2012_p2;
wire   [0:0] and_ln88_21_fu_1988_p2;
wire   [0:0] xor_ln88_27_fu_2018_p2;
wire   [0:0] xor_ln88_25_fu_2006_p2;
wire   [0:0] xor_ln88_28_fu_2024_p2;
wire   [0:0] and_ln91_5_fu_2054_p2;
wire   [0:0] xor_ln91_63_fu_2066_p2;
wire   [0:0] xor_ln91_62_fu_2060_p2;
wire   [0:0] and_ln90_16_fu_2042_p2;
wire   [0:0] and_ln90_15_fu_2036_p2;
wire   [0:0] xor_ln91_66_fu_2084_p2;
wire   [0:0] and_ln90_17_fu_2048_p2;
wire   [0:0] xor_ln91_67_fu_2090_p2;
wire   [0:0] xor_ln91_65_fu_2078_p2;
wire   [0:0] xor_ln91_68_fu_2096_p2;
wire   [0:0] xor_ln91_64_fu_2072_p2;
wire   [0:0] xor_ln91_11_fu_2102_p2;
wire   [0:0] xor_ln88_29_fu_2030_p2;
wire   [0:0] xor_ln87_29_fu_1976_p2;
wire   [0:0] xor_ln86_17_fu_1922_p2;
wire   [0:0] xor_ln54_2_fu_2126_p2;
wire   [0:0] xor_ln54_3_fu_2132_p2;
wire   [0:0] xor_ln53_1_fu_2120_p2;
wire   [3:0] res_44_fu_1810_p5;
wire   [3:0] res_43_fu_1496_p5;
wire   [3:0] res_45_fu_2108_p5;
wire   [3:0] res_4_fu_2138_p5;
wire   [3:0] xor_ln101_5_fu_2156_p2;
wire   [3:0] xor_ln101_4_fu_2150_p2;
wire   [3:0] xor_ln101_6_fu_2162_p2;
wire   [3:0] xor_ln101_7_fu_2168_p2;
wire   [0:0] tmp_40_fu_2202_p3;
wire   [0:0] tmp_41_fu_2210_p3;
wire   [0:0] tmp_42_fu_2224_p3;
wire   [0:0] tmp_43_fu_2232_p3;
wire   [0:0] tmp_44_fu_2246_p3;
wire   [0:0] tmp_45_fu_2254_p3;
wire   [0:0] tmp_46_fu_2268_p3;
wire   [0:0] tmp_47_fu_2276_p3;
wire   [0:0] and_ln86_24_fu_2218_p2;
wire   [0:0] and_ln86_25_fu_2240_p2;
wire   [0:0] and_ln86_26_fu_2262_p2;
wire   [0:0] and_ln86_27_fu_2284_p2;
wire   [0:0] xor_ln86_19_fu_2296_p2;
wire   [0:0] xor_ln86_18_fu_2290_p2;
wire   [0:0] and_ln87_25_fu_2314_p2;
wire   [0:0] xor_ln87_30_fu_2332_p2;
wire   [0:0] and_ln87_24_fu_2308_p2;
wire   [0:0] and_ln87_27_fu_2326_p2;
wire   [0:0] xor_ln87_32_fu_2344_p2;
wire   [0:0] and_ln87_26_fu_2320_p2;
wire   [0:0] xor_ln87_33_fu_2350_p2;
wire   [0:0] xor_ln87_31_fu_2338_p2;
wire   [0:0] and_ln88_25_fu_2368_p2;
wire   [0:0] and_ln88_26_fu_2374_p2;
wire   [0:0] xor_ln88_30_fu_2386_p2;
wire   [0:0] and_ln88_24_fu_2362_p2;
wire   [0:0] and_ln88_27_fu_2380_p2;
wire   [0:0] xor_ln88_32_fu_2398_p2;
wire   [0:0] xor_ln88_33_fu_2404_p2;
wire   [0:0] xor_ln88_31_fu_2392_p2;
wire   [0:0] and_ln90_18_fu_2416_p2;
wire   [0:0] and_ln90_19_fu_2422_p2;
wire   [0:0] and_ln90_20_fu_2428_p2;
wire   [0:0] xor_ln91_70_fu_2446_p2;
wire   [0:0] xor_ln91_69_fu_2440_p2;
wire   [0:0] xor_ln91_73_fu_2464_p2;
wire   [0:0] and_ln91_6_fu_2434_p2;
wire   [0:0] xor_ln91_74_fu_2470_p2;
wire   [0:0] xor_ln91_72_fu_2458_p2;
wire   [0:0] xor_ln91_75_fu_2476_p2;
wire   [0:0] xor_ln91_71_fu_2452_p2;
wire   [0:0] xor_ln91_13_fu_2482_p2;
wire   [0:0] xor_ln88_34_fu_2410_p2;
wire   [0:0] xor_ln87_34_fu_2356_p2;
wire   [0:0] xor_ln86_20_fu_2302_p2;
wire   [3:0] a1_14_fu_2182_p4;
wire   [3:0] b1_14_fu_2192_p4;
wire   [3:0] a_13_fu_2500_p2;
wire   [3:0] b_11_fu_2506_p2;
wire   [0:0] trunc_ln86_8_fu_2512_p1;
wire   [0:0] trunc_ln86_9_fu_2516_p1;
wire   [0:0] tmp_48_fu_2526_p3;
wire   [0:0] tmp_49_fu_2534_p3;
wire   [0:0] tmp_50_fu_2548_p3;
wire   [0:0] tmp_51_fu_2556_p3;
wire   [0:0] tmp_52_fu_2570_p3;
wire   [0:0] tmp_53_fu_2578_p3;
wire   [0:0] and_ln86_28_fu_2520_p2;
wire   [0:0] and_ln86_29_fu_2542_p2;
wire   [0:0] and_ln86_30_fu_2564_p2;
wire   [0:0] and_ln86_31_fu_2586_p2;
wire   [0:0] xor_ln86_22_fu_2598_p2;
wire   [0:0] xor_ln86_21_fu_2592_p2;
wire   [0:0] and_ln87_29_fu_2616_p2;
wire   [0:0] xor_ln87_35_fu_2634_p2;
wire   [0:0] and_ln87_28_fu_2610_p2;
wire   [0:0] and_ln87_31_fu_2628_p2;
wire   [0:0] xor_ln87_37_fu_2646_p2;
wire   [0:0] and_ln87_30_fu_2622_p2;
wire   [0:0] xor_ln87_38_fu_2652_p2;
wire   [0:0] xor_ln87_36_fu_2640_p2;
wire   [0:0] and_ln88_29_fu_2670_p2;
wire   [0:0] and_ln88_30_fu_2676_p2;
wire   [0:0] xor_ln88_35_fu_2688_p2;
wire   [0:0] and_ln88_28_fu_2664_p2;
wire   [0:0] and_ln88_31_fu_2682_p2;
wire   [0:0] xor_ln88_37_fu_2700_p2;
wire   [0:0] xor_ln88_38_fu_2706_p2;
wire   [0:0] xor_ln88_36_fu_2694_p2;
wire   [0:0] and_ln90_21_fu_2718_p2;
wire   [0:0] and_ln90_22_fu_2724_p2;
wire   [0:0] and_ln90_23_fu_2730_p2;
wire   [0:0] xor_ln91_77_fu_2748_p2;
wire   [0:0] xor_ln91_76_fu_2742_p2;
wire   [0:0] xor_ln91_80_fu_2766_p2;
wire   [0:0] and_ln91_7_fu_2736_p2;
wire   [0:0] xor_ln91_81_fu_2772_p2;
wire   [0:0] xor_ln91_79_fu_2760_p2;
wire   [0:0] xor_ln91_82_fu_2778_p2;
wire   [0:0] xor_ln91_78_fu_2754_p2;
wire   [0:0] xor_ln91_15_fu_2784_p2;
wire   [0:0] xor_ln88_39_fu_2712_p2;
wire   [0:0] xor_ln87_39_fu_2658_p2;
wire   [0:0] xor_ln86_23_fu_2604_p2;
wire   [0:0] tmp_54_fu_2802_p3;
wire   [0:0] tmp_55_fu_2810_p3;
wire   [0:0] tmp_56_fu_2824_p3;
wire   [0:0] tmp_57_fu_2832_p3;
wire   [0:0] tmp_58_fu_2846_p3;
wire   [0:0] tmp_59_fu_2854_p3;
wire   [0:0] tmp_60_fu_2868_p3;
wire   [0:0] tmp_61_fu_2876_p3;
wire   [0:0] and_ln86_33_fu_2840_p2;
wire   [0:0] and_ln86_34_fu_2862_p2;
wire   [0:0] and_ln86_32_fu_2818_p2;
wire   [0:0] and_ln86_35_fu_2884_p2;
wire   [0:0] xor_ln86_25_fu_2896_p2;
wire   [0:0] xor_ln86_24_fu_2890_p2;
wire   [0:0] and_ln87_33_fu_2914_p2;
wire   [0:0] and_ln87_32_fu_2908_p2;
wire   [0:0] and_ln87_34_fu_2920_p2;
wire   [0:0] xor_ln87_41_fu_2932_p2;
wire   [0:0] xor_ln87_40_fu_2926_p2;
wire   [0:0] and_ln87_35_fu_2944_p2;
wire   [0:0] xor_ln87_43_fu_2950_p2;
wire   [0:0] xor_ln87_42_fu_2938_p2;
wire   [0:0] and_ln88_34_fu_2974_p2;
wire   [0:0] and_ln88_32_fu_2962_p2;
wire   [0:0] and_ln88_35_fu_2980_p2;
wire   [0:0] xor_ln88_41_fu_2992_p2;
wire   [0:0] and_ln88_33_fu_2968_p2;
wire   [0:0] xor_ln88_42_fu_2998_p2;
wire   [0:0] xor_ln88_40_fu_2986_p2;
wire   [0:0] xor_ln88_43_fu_3004_p2;
wire   [0:0] and_ln91_8_fu_3034_p2;
wire   [0:0] xor_ln91_84_fu_3046_p2;
wire   [0:0] xor_ln91_83_fu_3040_p2;
wire   [0:0] and_ln90_25_fu_3022_p2;
wire   [0:0] and_ln90_24_fu_3016_p2;
wire   [0:0] xor_ln91_87_fu_3064_p2;
wire   [0:0] and_ln90_26_fu_3028_p2;
wire   [0:0] xor_ln91_88_fu_3070_p2;
wire   [0:0] xor_ln91_86_fu_3058_p2;
wire   [0:0] xor_ln91_89_fu_3076_p2;
wire   [0:0] xor_ln91_85_fu_3052_p2;
wire   [0:0] xor_ln91_17_fu_3082_p2;
wire   [0:0] xor_ln88_44_fu_3010_p2;
wire   [0:0] xor_ln87_44_fu_2956_p2;
wire   [0:0] xor_ln86_26_fu_2902_p2;
wire   [0:0] xor_ln54_4_fu_3106_p2;
wire   [0:0] xor_ln54_5_fu_3112_p2;
wire   [0:0] xor_ln53_2_fu_3100_p2;
wire   [3:0] res_46_fu_2488_p5;
wire   [3:0] res_48_fu_3088_p5;
wire   [3:0] res_47_fu_2790_p5;
wire   [3:0] res_8_fu_3118_p5;
wire   [3:0] xor_ln101_9_fu_3136_p2;
wire   [3:0] xor_ln101_8_fu_3130_p2;
wire   [3:0] xor_ln101_10_fu_3142_p2;
wire   [0:0] trunc_ln62_fu_3156_p1;
wire   [0:0] tmp_62_fu_3160_p3;
wire   [0:0] tmp_63_fu_3174_p3;
wire   [0:0] tmp_64_fu_3182_p3;
wire   [0:0] trunc_ln64_fu_3204_p1;
wire   [0:0] xor_ln64_fu_3208_p2;
wire   [0:0] tmp_65_fu_3196_p3;
wire   [0:0] tmp_66_fu_3220_p3;
wire   [0:0] tmp_67_fu_3228_p3;
wire   [0:0] xor_ln65_1_fu_3242_p2;
wire   [0:0] xor_ln65_fu_3236_p2;
wire   [0:0] xor_ln65_2_fu_3248_p2;
wire   [0:0] xor_ln64_1_fu_3214_p2;
wire   [0:0] xor_ln63_fu_3190_p2;
wire   [0:0] xor_ln62_fu_3168_p2;
wire   [7:0] z1_2_fu_2174_p3;
wire   [7:0] z0_1_fu_1158_p3;
wire   [7:0] z2_fu_3148_p3;
wire   [7:0] res_9_fu_3254_p6;
wire   [7:0] xor_ln101_12_fu_3274_p2;
wire   [7:0] xor_ln101_11_fu_3268_p2;
wire   [7:0] xor_ln101_13_fu_3280_p2;
wire   [7:0] xor_ln101_14_fu_3286_p2;
wire   [15:0] a1_fu_134_p4;
wire   [15:0] a0_11_fu_130_p1;
wire   [15:0] b1_fu_148_p4;
wire   [15:0] b0_fu_144_p1;
wire   [7:0] a0_18_fu_3310_p4;
wire   [15:0] a_17_fu_3320_p2;
wire   [7:0] b0_7_fu_3336_p4;
wire   [15:0] b_13_fu_3346_p2;
wire   [3:0] a0_19_fu_3300_p4;
wire   [7:0] a0_15_fu_3352_p2;
wire   [3:0] b0_8_fu_3326_p4;
wire   [7:0] b0_4_fu_3368_p2;
wire   [0:0] trunc_ln86_10_fu_3416_p1;
wire   [0:0] trunc_ln86_11_fu_3420_p1;
wire   [0:0] tmp_68_fu_3430_p3;
wire   [0:0] tmp_69_fu_3438_p3;
wire   [0:0] tmp_70_fu_3452_p3;
wire   [0:0] tmp_71_fu_3460_p3;
wire   [0:0] tmp_72_fu_3474_p3;
wire   [0:0] tmp_73_fu_3482_p3;
wire   [0:0] and_ln86_36_fu_3424_p2;
wire   [0:0] and_ln86_37_fu_3446_p2;
wire   [0:0] and_ln86_38_fu_3468_p2;
wire   [0:0] and_ln86_39_fu_3490_p2;
wire   [0:0] xor_ln86_28_fu_3502_p2;
wire   [0:0] xor_ln86_27_fu_3496_p2;
wire   [0:0] and_ln87_37_fu_3520_p2;
wire   [0:0] xor_ln87_45_fu_3538_p2;
wire   [0:0] and_ln87_36_fu_3514_p2;
wire   [0:0] and_ln87_39_fu_3532_p2;
wire   [0:0] xor_ln87_47_fu_3550_p2;
wire   [0:0] and_ln87_38_fu_3526_p2;
wire   [0:0] xor_ln87_48_fu_3556_p2;
wire   [0:0] xor_ln87_46_fu_3544_p2;
wire   [0:0] and_ln88_37_fu_3574_p2;
wire   [0:0] and_ln88_38_fu_3580_p2;
wire   [0:0] xor_ln88_45_fu_3592_p2;
wire   [0:0] and_ln88_36_fu_3568_p2;
wire   [0:0] and_ln88_39_fu_3586_p2;
wire   [0:0] xor_ln88_47_fu_3604_p2;
wire   [0:0] xor_ln88_48_fu_3610_p2;
wire   [0:0] xor_ln88_46_fu_3598_p2;
wire   [0:0] and_ln90_27_fu_3622_p2;
wire   [0:0] and_ln90_28_fu_3628_p2;
wire   [0:0] and_ln90_29_fu_3634_p2;
wire   [0:0] xor_ln91_91_fu_3652_p2;
wire   [0:0] xor_ln91_90_fu_3646_p2;
wire   [0:0] xor_ln91_94_fu_3670_p2;
wire   [0:0] and_ln91_9_fu_3640_p2;
wire   [0:0] xor_ln91_95_fu_3676_p2;
wire   [0:0] xor_ln91_93_fu_3664_p2;
wire   [0:0] xor_ln91_96_fu_3682_p2;
wire   [0:0] xor_ln91_92_fu_3658_p2;
wire   [0:0] xor_ln91_19_fu_3688_p2;
wire   [0:0] xor_ln88_49_fu_3616_p2;
wire   [0:0] xor_ln87_49_fu_3562_p2;
wire   [0:0] xor_ln86_29_fu_3508_p2;
wire   [3:0] a1_16_fu_3390_p4;
wire   [3:0] a0_16_fu_3384_p2;
wire   [3:0] b1_16_fu_3406_p4;
wire   [3:0] b0_5_fu_3400_p2;
wire   [3:0] a_20_fu_3706_p2;
wire   [3:0] b_16_fu_3712_p2;
wire   [0:0] trunc_ln86_12_fu_3718_p1;
wire   [0:0] trunc_ln86_13_fu_3722_p1;
wire   [0:0] tmp_74_fu_3732_p3;
wire   [0:0] tmp_75_fu_3740_p3;
wire   [0:0] tmp_76_fu_3754_p3;
wire   [0:0] tmp_77_fu_3762_p3;
wire   [0:0] tmp_78_fu_3776_p3;
wire   [0:0] tmp_79_fu_3784_p3;
wire   [0:0] and_ln86_40_fu_3726_p2;
wire   [0:0] and_ln86_41_fu_3748_p2;
wire   [0:0] and_ln86_42_fu_3770_p2;
wire   [0:0] and_ln86_43_fu_3792_p2;
wire   [0:0] xor_ln86_31_fu_3804_p2;
wire   [0:0] xor_ln86_30_fu_3798_p2;
wire   [0:0] and_ln87_41_fu_3822_p2;
wire   [0:0] xor_ln87_50_fu_3840_p2;
wire   [0:0] and_ln87_40_fu_3816_p2;
wire   [0:0] and_ln87_43_fu_3834_p2;
wire   [0:0] xor_ln87_52_fu_3852_p2;
wire   [0:0] and_ln87_42_fu_3828_p2;
wire   [0:0] xor_ln87_53_fu_3858_p2;
wire   [0:0] xor_ln87_51_fu_3846_p2;
wire   [0:0] and_ln88_41_fu_3876_p2;
wire   [0:0] and_ln88_42_fu_3882_p2;
wire   [0:0] xor_ln88_50_fu_3894_p2;
wire   [0:0] and_ln88_40_fu_3870_p2;
wire   [0:0] and_ln88_43_fu_3888_p2;
wire   [0:0] xor_ln88_52_fu_3906_p2;
wire   [0:0] xor_ln88_53_fu_3912_p2;
wire   [0:0] xor_ln88_51_fu_3900_p2;
wire   [0:0] and_ln90_30_fu_3924_p2;
wire   [0:0] and_ln90_31_fu_3930_p2;
wire   [0:0] and_ln90_32_fu_3936_p2;
wire   [0:0] xor_ln91_98_fu_3954_p2;
wire   [0:0] xor_ln91_97_fu_3948_p2;
wire   [0:0] xor_ln91_101_fu_3972_p2;
wire   [0:0] and_ln91_10_fu_3942_p2;
wire   [0:0] xor_ln91_102_fu_3978_p2;
wire   [0:0] xor_ln91_100_fu_3966_p2;
wire   [0:0] xor_ln91_103_fu_3984_p2;
wire   [0:0] xor_ln91_99_fu_3960_p2;
wire   [0:0] xor_ln91_21_fu_3990_p2;
wire   [0:0] xor_ln88_54_fu_3918_p2;
wire   [0:0] xor_ln87_54_fu_3864_p2;
wire   [0:0] xor_ln86_32_fu_3810_p2;
wire   [0:0] tmp_80_fu_4008_p3;
wire   [0:0] tmp_81_fu_4016_p3;
wire   [0:0] tmp_82_fu_4030_p3;
wire   [0:0] tmp_83_fu_4038_p3;
wire   [0:0] tmp_84_fu_4052_p3;
wire   [0:0] tmp_85_fu_4060_p3;
wire   [0:0] tmp_86_fu_4074_p3;
wire   [0:0] tmp_87_fu_4082_p3;
wire   [0:0] and_ln86_45_fu_4046_p2;
wire   [0:0] and_ln86_46_fu_4068_p2;
wire   [0:0] and_ln86_44_fu_4024_p2;
wire   [0:0] and_ln86_47_fu_4090_p2;
wire   [0:0] xor_ln86_34_fu_4102_p2;
wire   [0:0] xor_ln86_33_fu_4096_p2;
wire   [0:0] and_ln87_45_fu_4120_p2;
wire   [0:0] and_ln87_44_fu_4114_p2;
wire   [0:0] and_ln87_46_fu_4126_p2;
wire   [0:0] xor_ln87_56_fu_4138_p2;
wire   [0:0] xor_ln87_55_fu_4132_p2;
wire   [0:0] and_ln87_47_fu_4150_p2;
wire   [0:0] xor_ln87_58_fu_4156_p2;
wire   [0:0] xor_ln87_57_fu_4144_p2;
wire   [0:0] and_ln88_46_fu_4180_p2;
wire   [0:0] and_ln88_44_fu_4168_p2;
wire   [0:0] and_ln88_47_fu_4186_p2;
wire   [0:0] xor_ln88_56_fu_4198_p2;
wire   [0:0] and_ln88_45_fu_4174_p2;
wire   [0:0] xor_ln88_57_fu_4204_p2;
wire   [0:0] xor_ln88_55_fu_4192_p2;
wire   [0:0] xor_ln88_58_fu_4210_p2;
wire   [0:0] and_ln91_11_fu_4240_p2;
wire   [0:0] xor_ln91_105_fu_4252_p2;
wire   [0:0] xor_ln91_104_fu_4246_p2;
wire   [0:0] and_ln90_34_fu_4228_p2;
wire   [0:0] and_ln90_33_fu_4222_p2;
wire   [0:0] xor_ln91_108_fu_4270_p2;
wire   [0:0] and_ln90_35_fu_4234_p2;
wire   [0:0] xor_ln91_109_fu_4276_p2;
wire   [0:0] xor_ln91_107_fu_4264_p2;
wire   [0:0] xor_ln91_110_fu_4282_p2;
wire   [0:0] xor_ln91_106_fu_4258_p2;
wire   [0:0] xor_ln91_23_fu_4288_p2;
wire   [0:0] xor_ln88_59_fu_4216_p2;
wire   [0:0] xor_ln87_59_fu_4162_p2;
wire   [0:0] xor_ln86_35_fu_4108_p2;
wire   [0:0] xor_ln54_6_fu_4312_p2;
wire   [0:0] xor_ln54_7_fu_4318_p2;
wire   [0:0] xor_ln53_3_fu_4306_p2;
wire   [3:0] res_50_fu_3996_p5;
wire   [3:0] res_49_fu_3694_p5;
wire   [3:0] res_51_fu_4294_p5;
wire   [3:0] res_16_fu_4324_p5;
wire   [3:0] xor_ln101_16_fu_4342_p2;
wire   [3:0] xor_ln101_15_fu_4336_p2;
wire   [3:0] xor_ln101_17_fu_4348_p2;
wire   [3:0] xor_ln101_18_fu_4354_p2;
wire   [7:0] a1_15_fu_3358_p4;
wire   [7:0] b1_15_fu_3374_p4;
wire   [7:0] a_23_fu_4378_p2;
wire   [7:0] b_18_fu_4394_p2;
wire   [0:0] trunc_ln86_14_fu_4420_p1;
wire   [0:0] trunc_ln86_15_fu_4424_p1;
wire   [0:0] tmp_88_fu_4434_p3;
wire   [0:0] tmp_89_fu_4442_p3;
wire   [0:0] tmp_90_fu_4456_p3;
wire   [0:0] tmp_91_fu_4464_p3;
wire   [0:0] tmp_92_fu_4478_p3;
wire   [0:0] tmp_93_fu_4486_p3;
wire   [0:0] and_ln86_48_fu_4428_p2;
wire   [0:0] and_ln86_49_fu_4450_p2;
wire   [0:0] and_ln86_50_fu_4472_p2;
wire   [0:0] and_ln86_51_fu_4494_p2;
wire   [0:0] xor_ln86_37_fu_4506_p2;
wire   [0:0] xor_ln86_36_fu_4500_p2;
wire   [0:0] and_ln87_49_fu_4524_p2;
wire   [0:0] xor_ln87_60_fu_4542_p2;
wire   [0:0] and_ln87_48_fu_4518_p2;
wire   [0:0] and_ln87_51_fu_4536_p2;
wire   [0:0] xor_ln87_62_fu_4554_p2;
wire   [0:0] and_ln87_50_fu_4530_p2;
wire   [0:0] xor_ln87_63_fu_4560_p2;
wire   [0:0] xor_ln87_61_fu_4548_p2;
wire   [0:0] and_ln88_49_fu_4578_p2;
wire   [0:0] and_ln88_50_fu_4584_p2;
wire   [0:0] xor_ln88_60_fu_4596_p2;
wire   [0:0] and_ln88_48_fu_4572_p2;
wire   [0:0] and_ln88_51_fu_4590_p2;
wire   [0:0] xor_ln88_62_fu_4608_p2;
wire   [0:0] xor_ln88_63_fu_4614_p2;
wire   [0:0] xor_ln88_61_fu_4602_p2;
wire   [0:0] and_ln90_36_fu_4626_p2;
wire   [0:0] and_ln90_37_fu_4632_p2;
wire   [0:0] and_ln90_38_fu_4638_p2;
wire   [0:0] xor_ln91_112_fu_4656_p2;
wire   [0:0] xor_ln91_111_fu_4650_p2;
wire   [0:0] xor_ln91_115_fu_4674_p2;
wire   [0:0] and_ln91_12_fu_4644_p2;
wire   [0:0] xor_ln91_116_fu_4680_p2;
wire   [0:0] xor_ln91_114_fu_4668_p2;
wire   [0:0] xor_ln91_117_fu_4686_p2;
wire   [0:0] xor_ln91_113_fu_4662_p2;
wire   [0:0] xor_ln91_25_fu_4692_p2;
wire   [0:0] xor_ln88_64_fu_4620_p2;
wire   [0:0] xor_ln87_64_fu_4566_p2;
wire   [0:0] xor_ln86_38_fu_4512_p2;
wire   [3:0] a1_17_fu_4400_p4;
wire   [3:0] xor_ln99_14_fu_4710_p2;
wire   [3:0] a0_17_fu_4368_p4;
wire   [3:0] b1_17_fu_4410_p4;
wire   [3:0] xor_ln99_16_fu_4722_p2;
wire   [3:0] b0_6_fu_4384_p4;
wire   [3:0] a_24_fu_4716_p2;
wire   [3:0] b_19_fu_4728_p2;
wire   [0:0] trunc_ln86_16_fu_4734_p1;
wire   [0:0] trunc_ln86_17_fu_4738_p1;
wire   [0:0] tmp_94_fu_4748_p3;
wire   [0:0] tmp_95_fu_4756_p3;
wire   [0:0] tmp_96_fu_4770_p3;
wire   [0:0] tmp_97_fu_4778_p3;
wire   [0:0] tmp_98_fu_4792_p3;
wire   [0:0] tmp_99_fu_4800_p3;
wire   [0:0] and_ln86_52_fu_4742_p2;
wire   [0:0] and_ln86_53_fu_4764_p2;
wire   [0:0] and_ln86_54_fu_4786_p2;
wire   [0:0] and_ln86_55_fu_4808_p2;
wire   [0:0] xor_ln86_40_fu_4820_p2;
wire   [0:0] xor_ln86_39_fu_4814_p2;
wire   [0:0] and_ln87_53_fu_4838_p2;
wire   [0:0] xor_ln87_65_fu_4856_p2;
wire   [0:0] and_ln87_52_fu_4832_p2;
wire   [0:0] and_ln87_55_fu_4850_p2;
wire   [0:0] xor_ln87_67_fu_4868_p2;
wire   [0:0] and_ln87_54_fu_4844_p2;
wire   [0:0] xor_ln87_68_fu_4874_p2;
wire   [0:0] xor_ln87_66_fu_4862_p2;
wire   [0:0] and_ln88_53_fu_4892_p2;
wire   [0:0] and_ln88_54_fu_4898_p2;
wire   [0:0] xor_ln88_65_fu_4910_p2;
wire   [0:0] and_ln88_52_fu_4886_p2;
wire   [0:0] and_ln88_55_fu_4904_p2;
wire   [0:0] xor_ln88_67_fu_4922_p2;
wire   [0:0] xor_ln88_68_fu_4928_p2;
wire   [0:0] xor_ln88_66_fu_4916_p2;
wire   [0:0] and_ln90_39_fu_4940_p2;
wire   [0:0] and_ln90_40_fu_4946_p2;
wire   [0:0] and_ln90_41_fu_4952_p2;
wire   [0:0] xor_ln91_119_fu_4970_p2;
wire   [0:0] xor_ln91_118_fu_4964_p2;
wire   [0:0] xor_ln91_122_fu_4988_p2;
wire   [0:0] and_ln91_13_fu_4958_p2;
wire   [0:0] xor_ln91_123_fu_4994_p2;
wire   [0:0] xor_ln91_121_fu_4982_p2;
wire   [0:0] xor_ln91_124_fu_5000_p2;
wire   [0:0] xor_ln91_120_fu_4976_p2;
wire   [0:0] xor_ln91_27_fu_5006_p2;
wire   [0:0] xor_ln88_69_fu_4934_p2;
wire   [0:0] xor_ln87_69_fu_4880_p2;
wire   [0:0] xor_ln86_41_fu_4826_p2;
wire   [0:0] tmp_100_fu_5024_p3;
wire   [0:0] tmp_101_fu_5032_p3;
wire   [0:0] tmp_102_fu_5046_p3;
wire   [0:0] tmp_103_fu_5054_p3;
wire   [0:0] tmp_104_fu_5068_p3;
wire   [0:0] tmp_105_fu_5076_p3;
wire   [0:0] tmp_106_fu_5090_p3;
wire   [0:0] tmp_107_fu_5098_p3;
wire   [0:0] and_ln86_57_fu_5062_p2;
wire   [0:0] and_ln86_58_fu_5084_p2;
wire   [0:0] and_ln86_56_fu_5040_p2;
wire   [0:0] and_ln86_59_fu_5106_p2;
wire   [0:0] xor_ln86_43_fu_5118_p2;
wire   [0:0] xor_ln86_42_fu_5112_p2;
wire   [0:0] and_ln87_57_fu_5136_p2;
wire   [0:0] and_ln87_56_fu_5130_p2;
wire   [0:0] and_ln87_58_fu_5142_p2;
wire   [0:0] xor_ln87_71_fu_5154_p2;
wire   [0:0] xor_ln87_70_fu_5148_p2;
wire   [0:0] and_ln87_59_fu_5166_p2;
wire   [0:0] xor_ln87_73_fu_5172_p2;
wire   [0:0] xor_ln87_72_fu_5160_p2;
wire   [0:0] and_ln88_58_fu_5196_p2;
wire   [0:0] and_ln88_56_fu_5184_p2;
wire   [0:0] and_ln88_59_fu_5202_p2;
wire   [0:0] xor_ln88_71_fu_5214_p2;
wire   [0:0] and_ln88_57_fu_5190_p2;
wire   [0:0] xor_ln88_72_fu_5220_p2;
wire   [0:0] xor_ln88_70_fu_5208_p2;
wire   [0:0] xor_ln88_73_fu_5226_p2;
wire   [0:0] and_ln91_14_fu_5256_p2;
wire   [0:0] xor_ln91_126_fu_5268_p2;
wire   [0:0] xor_ln91_125_fu_5262_p2;
wire   [0:0] and_ln90_43_fu_5244_p2;
wire   [0:0] and_ln90_42_fu_5238_p2;
wire   [0:0] xor_ln91_129_fu_5286_p2;
wire   [0:0] and_ln90_44_fu_5250_p2;
wire   [0:0] xor_ln91_130_fu_5292_p2;
wire   [0:0] xor_ln91_128_fu_5280_p2;
wire   [0:0] xor_ln91_131_fu_5298_p2;
wire   [0:0] xor_ln91_127_fu_5274_p2;
wire   [0:0] xor_ln91_29_fu_5304_p2;
wire   [0:0] xor_ln88_74_fu_5232_p2;
wire   [0:0] xor_ln87_74_fu_5178_p2;
wire   [0:0] xor_ln86_44_fu_5124_p2;
wire   [0:0] xor_ln54_8_fu_5328_p2;
wire   [0:0] xor_ln54_9_fu_5334_p2;
wire   [0:0] xor_ln53_4_fu_5322_p2;
wire   [3:0] res_53_fu_5012_p5;
wire   [3:0] res_52_fu_4698_p5;
wire   [3:0] res_54_fu_5310_p5;
wire   [3:0] res_20_fu_5340_p5;
wire   [3:0] xor_ln101_20_fu_5358_p2;
wire   [3:0] xor_ln101_19_fu_5352_p2;
wire   [3:0] xor_ln101_21_fu_5364_p2;
wire   [3:0] xor_ln101_22_fu_5370_p2;
wire   [0:0] tmp_108_fu_5404_p3;
wire   [0:0] tmp_109_fu_5412_p3;
wire   [0:0] tmp_110_fu_5426_p3;
wire   [0:0] tmp_111_fu_5434_p3;
wire   [0:0] tmp_112_fu_5448_p3;
wire   [0:0] tmp_113_fu_5456_p3;
wire   [0:0] tmp_114_fu_5470_p3;
wire   [0:0] tmp_115_fu_5478_p3;
wire   [0:0] and_ln86_60_fu_5420_p2;
wire   [0:0] and_ln86_61_fu_5442_p2;
wire   [0:0] and_ln86_62_fu_5464_p2;
wire   [0:0] and_ln86_63_fu_5486_p2;
wire   [0:0] xor_ln86_46_fu_5498_p2;
wire   [0:0] xor_ln86_45_fu_5492_p2;
wire   [0:0] and_ln87_61_fu_5516_p2;
wire   [0:0] xor_ln87_75_fu_5534_p2;
wire   [0:0] and_ln87_60_fu_5510_p2;
wire   [0:0] and_ln87_63_fu_5528_p2;
wire   [0:0] xor_ln87_77_fu_5546_p2;
wire   [0:0] and_ln87_62_fu_5522_p2;
wire   [0:0] xor_ln87_78_fu_5552_p2;
wire   [0:0] xor_ln87_76_fu_5540_p2;
wire   [0:0] and_ln88_61_fu_5570_p2;
wire   [0:0] and_ln88_62_fu_5576_p2;
wire   [0:0] xor_ln88_75_fu_5588_p2;
wire   [0:0] and_ln88_60_fu_5564_p2;
wire   [0:0] and_ln88_63_fu_5582_p2;
wire   [0:0] xor_ln88_77_fu_5600_p2;
wire   [0:0] xor_ln88_78_fu_5606_p2;
wire   [0:0] xor_ln88_76_fu_5594_p2;
wire   [0:0] and_ln90_45_fu_5618_p2;
wire   [0:0] and_ln90_46_fu_5624_p2;
wire   [0:0] and_ln90_47_fu_5630_p2;
wire   [0:0] xor_ln91_133_fu_5648_p2;
wire   [0:0] xor_ln91_132_fu_5642_p2;
wire   [0:0] xor_ln91_136_fu_5666_p2;
wire   [0:0] and_ln91_15_fu_5636_p2;
wire   [0:0] xor_ln91_137_fu_5672_p2;
wire   [0:0] xor_ln91_135_fu_5660_p2;
wire   [0:0] xor_ln91_138_fu_5678_p2;
wire   [0:0] xor_ln91_134_fu_5654_p2;
wire   [0:0] xor_ln91_31_fu_5684_p2;
wire   [0:0] xor_ln88_79_fu_5612_p2;
wire   [0:0] xor_ln87_79_fu_5558_p2;
wire   [0:0] xor_ln86_47_fu_5504_p2;
wire   [3:0] a1_18_fu_5384_p4;
wire   [3:0] b1_18_fu_5394_p4;
wire   [3:0] a_29_fu_5702_p2;
wire   [3:0] b_23_fu_5708_p2;
wire   [0:0] trunc_ln86_18_fu_5714_p1;
wire   [0:0] trunc_ln86_19_fu_5718_p1;
wire   [0:0] tmp_116_fu_5728_p3;
wire   [0:0] tmp_117_fu_5736_p3;
wire   [0:0] tmp_118_fu_5750_p3;
wire   [0:0] tmp_119_fu_5758_p3;
wire   [0:0] tmp_120_fu_5772_p3;
wire   [0:0] tmp_121_fu_5780_p3;
wire   [0:0] and_ln86_64_fu_5722_p2;
wire   [0:0] and_ln86_65_fu_5744_p2;
wire   [0:0] and_ln86_66_fu_5766_p2;
wire   [0:0] and_ln86_67_fu_5788_p2;
wire   [0:0] xor_ln86_49_fu_5800_p2;
wire   [0:0] xor_ln86_48_fu_5794_p2;
wire   [0:0] and_ln87_65_fu_5818_p2;
wire   [0:0] xor_ln87_80_fu_5836_p2;
wire   [0:0] and_ln87_64_fu_5812_p2;
wire   [0:0] and_ln87_67_fu_5830_p2;
wire   [0:0] xor_ln87_82_fu_5848_p2;
wire   [0:0] and_ln87_66_fu_5824_p2;
wire   [0:0] xor_ln87_83_fu_5854_p2;
wire   [0:0] xor_ln87_81_fu_5842_p2;
wire   [0:0] and_ln88_65_fu_5872_p2;
wire   [0:0] and_ln88_66_fu_5878_p2;
wire   [0:0] xor_ln88_80_fu_5890_p2;
wire   [0:0] and_ln88_64_fu_5866_p2;
wire   [0:0] and_ln88_67_fu_5884_p2;
wire   [0:0] xor_ln88_82_fu_5902_p2;
wire   [0:0] xor_ln88_83_fu_5908_p2;
wire   [0:0] xor_ln88_81_fu_5896_p2;
wire   [0:0] and_ln90_48_fu_5920_p2;
wire   [0:0] and_ln90_49_fu_5926_p2;
wire   [0:0] and_ln90_50_fu_5932_p2;
wire   [0:0] xor_ln91_140_fu_5950_p2;
wire   [0:0] xor_ln91_139_fu_5944_p2;
wire   [0:0] xor_ln91_143_fu_5968_p2;
wire   [0:0] and_ln91_16_fu_5938_p2;
wire   [0:0] xor_ln91_144_fu_5974_p2;
wire   [0:0] xor_ln91_142_fu_5962_p2;
wire   [0:0] xor_ln91_145_fu_5980_p2;
wire   [0:0] xor_ln91_141_fu_5956_p2;
wire   [0:0] xor_ln91_33_fu_5986_p2;
wire   [0:0] xor_ln88_84_fu_5914_p2;
wire   [0:0] xor_ln87_84_fu_5860_p2;
wire   [0:0] xor_ln86_50_fu_5806_p2;
wire   [0:0] tmp_122_fu_6004_p3;
wire   [0:0] tmp_123_fu_6012_p3;
wire   [0:0] tmp_124_fu_6026_p3;
wire   [0:0] tmp_125_fu_6034_p3;
wire   [0:0] tmp_126_fu_6048_p3;
wire   [0:0] tmp_127_fu_6056_p3;
wire   [0:0] tmp_128_fu_6070_p3;
wire   [0:0] tmp_129_fu_6078_p3;
wire   [0:0] and_ln86_69_fu_6042_p2;
wire   [0:0] and_ln86_70_fu_6064_p2;
wire   [0:0] and_ln86_68_fu_6020_p2;
wire   [0:0] and_ln86_71_fu_6086_p2;
wire   [0:0] xor_ln86_52_fu_6098_p2;
wire   [0:0] xor_ln86_51_fu_6092_p2;
wire   [0:0] and_ln87_69_fu_6116_p2;
wire   [0:0] and_ln87_68_fu_6110_p2;
wire   [0:0] and_ln87_70_fu_6122_p2;
wire   [0:0] xor_ln87_86_fu_6134_p2;
wire   [0:0] xor_ln87_85_fu_6128_p2;
wire   [0:0] and_ln87_71_fu_6146_p2;
wire   [0:0] xor_ln87_88_fu_6152_p2;
wire   [0:0] xor_ln87_87_fu_6140_p2;
wire   [0:0] and_ln88_70_fu_6176_p2;
wire   [0:0] and_ln88_68_fu_6164_p2;
wire   [0:0] and_ln88_71_fu_6182_p2;
wire   [0:0] xor_ln88_86_fu_6194_p2;
wire   [0:0] and_ln88_69_fu_6170_p2;
wire   [0:0] xor_ln88_87_fu_6200_p2;
wire   [0:0] xor_ln88_85_fu_6188_p2;
wire   [0:0] xor_ln88_88_fu_6206_p2;
wire   [0:0] and_ln91_17_fu_6236_p2;
wire   [0:0] xor_ln91_147_fu_6248_p2;
wire   [0:0] xor_ln91_146_fu_6242_p2;
wire   [0:0] and_ln90_52_fu_6224_p2;
wire   [0:0] and_ln90_51_fu_6218_p2;
wire   [0:0] xor_ln91_150_fu_6266_p2;
wire   [0:0] and_ln90_53_fu_6230_p2;
wire   [0:0] xor_ln91_151_fu_6272_p2;
wire   [0:0] xor_ln91_149_fu_6260_p2;
wire   [0:0] xor_ln91_152_fu_6278_p2;
wire   [0:0] xor_ln91_148_fu_6254_p2;
wire   [0:0] xor_ln91_35_fu_6284_p2;
wire   [0:0] xor_ln88_89_fu_6212_p2;
wire   [0:0] xor_ln87_89_fu_6158_p2;
wire   [0:0] xor_ln86_53_fu_6104_p2;
wire   [0:0] xor_ln54_10_fu_6308_p2;
wire   [0:0] xor_ln54_11_fu_6314_p2;
wire   [0:0] xor_ln53_5_fu_6302_p2;
wire   [3:0] res_55_fu_5690_p5;
wire   [3:0] res_57_fu_6290_p5;
wire   [3:0] res_56_fu_5992_p5;
wire   [3:0] res_24_fu_6320_p5;
wire   [3:0] xor_ln101_24_fu_6338_p2;
wire   [3:0] xor_ln101_23_fu_6332_p2;
wire   [3:0] xor_ln101_25_fu_6344_p2;
wire   [0:0] trunc_ln62_1_fu_6358_p1;
wire   [0:0] tmp_130_fu_6362_p3;
wire   [0:0] tmp_131_fu_6376_p3;
wire   [0:0] tmp_132_fu_6384_p3;
wire   [0:0] trunc_ln64_1_fu_6406_p1;
wire   [0:0] xor_ln64_2_fu_6410_p2;
wire   [0:0] tmp_133_fu_6398_p3;
wire   [0:0] tmp_134_fu_6422_p3;
wire   [0:0] tmp_135_fu_6430_p3;
wire   [0:0] xor_ln65_4_fu_6444_p2;
wire   [0:0] xor_ln65_3_fu_6438_p2;
wire   [0:0] xor_ln65_5_fu_6450_p2;
wire   [0:0] xor_ln64_3_fu_6416_p2;
wire   [0:0] xor_ln63_1_fu_6392_p2;
wire   [0:0] xor_ln62_1_fu_6370_p2;
wire   [7:0] z1_6_fu_5376_p3;
wire   [7:0] z0_6_fu_4360_p3;
wire   [7:0] z2_4_fu_6350_p3;
wire   [7:0] res_25_fu_6456_p6;
wire   [7:0] xor_ln101_27_fu_6476_p2;
wire   [7:0] xor_ln101_26_fu_6470_p2;
wire   [7:0] xor_ln101_28_fu_6482_p2;
wire   [7:0] xor_ln101_29_fu_6488_p2;
wire   [0:0] tmp_136_fu_6542_p3;
wire   [0:0] tmp_137_fu_6550_p3;
wire   [0:0] tmp_138_fu_6564_p3;
wire   [0:0] tmp_139_fu_6572_p3;
wire   [0:0] tmp_140_fu_6586_p3;
wire   [0:0] tmp_141_fu_6594_p3;
wire   [0:0] tmp_142_fu_6608_p3;
wire   [0:0] tmp_143_fu_6616_p3;
wire   [0:0] and_ln86_72_fu_6558_p2;
wire   [0:0] and_ln86_73_fu_6580_p2;
wire   [0:0] and_ln86_74_fu_6602_p2;
wire   [0:0] and_ln86_75_fu_6624_p2;
wire   [0:0] xor_ln86_55_fu_6636_p2;
wire   [0:0] xor_ln86_54_fu_6630_p2;
wire   [0:0] and_ln87_73_fu_6654_p2;
wire   [0:0] xor_ln87_90_fu_6672_p2;
wire   [0:0] and_ln87_72_fu_6648_p2;
wire   [0:0] and_ln87_75_fu_6666_p2;
wire   [0:0] xor_ln87_92_fu_6684_p2;
wire   [0:0] and_ln87_74_fu_6660_p2;
wire   [0:0] xor_ln87_93_fu_6690_p2;
wire   [0:0] xor_ln87_91_fu_6678_p2;
wire   [0:0] and_ln88_73_fu_6708_p2;
wire   [0:0] and_ln88_74_fu_6714_p2;
wire   [0:0] xor_ln88_90_fu_6726_p2;
wire   [0:0] and_ln88_72_fu_6702_p2;
wire   [0:0] and_ln88_75_fu_6720_p2;
wire   [0:0] xor_ln88_92_fu_6738_p2;
wire   [0:0] xor_ln88_93_fu_6744_p2;
wire   [0:0] xor_ln88_91_fu_6732_p2;
wire   [0:0] and_ln90_54_fu_6756_p2;
wire   [0:0] and_ln90_55_fu_6762_p2;
wire   [0:0] and_ln90_56_fu_6768_p2;
wire   [0:0] xor_ln91_154_fu_6786_p2;
wire   [0:0] xor_ln91_153_fu_6780_p2;
wire   [0:0] xor_ln91_157_fu_6804_p2;
wire   [0:0] and_ln91_18_fu_6774_p2;
wire   [0:0] xor_ln91_158_fu_6810_p2;
wire   [0:0] xor_ln91_156_fu_6798_p2;
wire   [0:0] xor_ln91_159_fu_6816_p2;
wire   [0:0] xor_ln91_155_fu_6792_p2;
wire   [0:0] xor_ln91_37_fu_6822_p2;
wire   [0:0] xor_ln88_94_fu_6750_p2;
wire   [0:0] xor_ln87_94_fu_6696_p2;
wire   [0:0] xor_ln86_56_fu_6642_p2;
wire   [3:0] a1_20_fu_6522_p4;
wire   [3:0] b1_20_fu_6532_p4;
wire   [3:0] a_36_fu_6840_p2;
wire   [3:0] b_28_fu_6846_p2;
wire   [0:0] trunc_ln86_20_fu_6852_p1;
wire   [0:0] trunc_ln86_21_fu_6856_p1;
wire   [0:0] tmp_144_fu_6866_p3;
wire   [0:0] tmp_145_fu_6874_p3;
wire   [0:0] tmp_146_fu_6888_p3;
wire   [0:0] tmp_147_fu_6896_p3;
wire   [0:0] tmp_148_fu_6910_p3;
wire   [0:0] tmp_149_fu_6918_p3;
wire   [0:0] and_ln86_76_fu_6860_p2;
wire   [0:0] and_ln86_77_fu_6882_p2;
wire   [0:0] and_ln86_78_fu_6904_p2;
wire   [0:0] and_ln86_79_fu_6926_p2;
wire   [0:0] xor_ln86_58_fu_6938_p2;
wire   [0:0] xor_ln86_57_fu_6932_p2;
wire   [0:0] and_ln87_77_fu_6956_p2;
wire   [0:0] xor_ln87_95_fu_6974_p2;
wire   [0:0] and_ln87_76_fu_6950_p2;
wire   [0:0] and_ln87_79_fu_6968_p2;
wire   [0:0] xor_ln87_97_fu_6986_p2;
wire   [0:0] and_ln87_78_fu_6962_p2;
wire   [0:0] xor_ln87_98_fu_6992_p2;
wire   [0:0] xor_ln87_96_fu_6980_p2;
wire   [0:0] and_ln88_77_fu_7010_p2;
wire   [0:0] and_ln88_78_fu_7016_p2;
wire   [0:0] xor_ln88_95_fu_7028_p2;
wire   [0:0] and_ln88_76_fu_7004_p2;
wire   [0:0] and_ln88_79_fu_7022_p2;
wire   [0:0] xor_ln88_97_fu_7040_p2;
wire   [0:0] xor_ln88_98_fu_7046_p2;
wire   [0:0] xor_ln88_96_fu_7034_p2;
wire   [0:0] and_ln90_57_fu_7058_p2;
wire   [0:0] and_ln90_58_fu_7064_p2;
wire   [0:0] and_ln90_59_fu_7070_p2;
wire   [0:0] xor_ln91_161_fu_7088_p2;
wire   [0:0] xor_ln91_160_fu_7082_p2;
wire   [0:0] xor_ln91_164_fu_7106_p2;
wire   [0:0] and_ln91_19_fu_7076_p2;
wire   [0:0] xor_ln91_165_fu_7112_p2;
wire   [0:0] xor_ln91_163_fu_7100_p2;
wire   [0:0] xor_ln91_166_fu_7118_p2;
wire   [0:0] xor_ln91_162_fu_7094_p2;
wire   [0:0] xor_ln91_39_fu_7124_p2;
wire   [0:0] xor_ln88_99_fu_7052_p2;
wire   [0:0] xor_ln87_99_fu_6998_p2;
wire   [0:0] xor_ln86_59_fu_6944_p2;
wire   [0:0] tmp_150_fu_7142_p3;
wire   [0:0] tmp_151_fu_7150_p3;
wire   [0:0] tmp_152_fu_7164_p3;
wire   [0:0] tmp_153_fu_7172_p3;
wire   [0:0] tmp_154_fu_7186_p3;
wire   [0:0] tmp_155_fu_7194_p3;
wire   [0:0] tmp_156_fu_7208_p3;
wire   [0:0] tmp_157_fu_7216_p3;
wire   [0:0] and_ln86_81_fu_7180_p2;
wire   [0:0] and_ln86_82_fu_7202_p2;
wire   [0:0] and_ln86_80_fu_7158_p2;
wire   [0:0] and_ln86_83_fu_7224_p2;
wire   [0:0] xor_ln86_61_fu_7236_p2;
wire   [0:0] xor_ln86_60_fu_7230_p2;
wire   [0:0] and_ln87_81_fu_7254_p2;
wire   [0:0] and_ln87_80_fu_7248_p2;
wire   [0:0] and_ln87_82_fu_7260_p2;
wire   [0:0] xor_ln87_101_fu_7272_p2;
wire   [0:0] xor_ln87_100_fu_7266_p2;
wire   [0:0] and_ln87_83_fu_7284_p2;
wire   [0:0] xor_ln87_103_fu_7290_p2;
wire   [0:0] xor_ln87_102_fu_7278_p2;
wire   [0:0] and_ln88_82_fu_7314_p2;
wire   [0:0] and_ln88_80_fu_7302_p2;
wire   [0:0] and_ln88_83_fu_7320_p2;
wire   [0:0] xor_ln88_101_fu_7332_p2;
wire   [0:0] and_ln88_81_fu_7308_p2;
wire   [0:0] xor_ln88_102_fu_7338_p2;
wire   [0:0] xor_ln88_100_fu_7326_p2;
wire   [0:0] xor_ln88_103_fu_7344_p2;
wire   [0:0] and_ln91_20_fu_7374_p2;
wire   [0:0] xor_ln91_168_fu_7386_p2;
wire   [0:0] xor_ln91_167_fu_7380_p2;
wire   [0:0] and_ln90_61_fu_7362_p2;
wire   [0:0] and_ln90_60_fu_7356_p2;
wire   [0:0] xor_ln91_171_fu_7404_p2;
wire   [0:0] and_ln90_62_fu_7368_p2;
wire   [0:0] xor_ln91_172_fu_7410_p2;
wire   [0:0] xor_ln91_170_fu_7398_p2;
wire   [0:0] xor_ln91_173_fu_7416_p2;
wire   [0:0] xor_ln91_169_fu_7392_p2;
wire   [0:0] xor_ln91_41_fu_7422_p2;
wire   [0:0] xor_ln88_104_fu_7350_p2;
wire   [0:0] xor_ln87_104_fu_7296_p2;
wire   [0:0] xor_ln86_62_fu_7242_p2;
wire   [0:0] xor_ln54_12_fu_7446_p2;
wire   [0:0] xor_ln54_13_fu_7452_p2;
wire   [0:0] xor_ln53_6_fu_7440_p2;
wire   [3:0] res_59_fu_7130_p5;
wire   [3:0] res_58_fu_6828_p5;
wire   [3:0] res_60_fu_7428_p5;
wire   [3:0] res_29_fu_7458_p5;
wire   [3:0] xor_ln101_31_fu_7476_p2;
wire   [3:0] xor_ln101_30_fu_7470_p2;
wire   [3:0] xor_ln101_32_fu_7482_p2;
wire   [3:0] xor_ln101_33_fu_7488_p2;
wire   [7:0] a1_19_fu_6502_p4;
wire   [7:0] b1_19_fu_6512_p4;
wire   [7:0] a_39_fu_7512_p2;
wire   [7:0] b_30_fu_7528_p2;
wire   [0:0] trunc_ln86_22_fu_7554_p1;
wire   [0:0] trunc_ln86_23_fu_7558_p1;
wire   [0:0] tmp_158_fu_7568_p3;
wire   [0:0] tmp_159_fu_7576_p3;
wire   [0:0] tmp_160_fu_7590_p3;
wire   [0:0] tmp_161_fu_7598_p3;
wire   [0:0] tmp_162_fu_7612_p3;
wire   [0:0] tmp_163_fu_7620_p3;
wire   [0:0] and_ln86_84_fu_7562_p2;
wire   [0:0] and_ln86_85_fu_7584_p2;
wire   [0:0] and_ln86_86_fu_7606_p2;
wire   [0:0] and_ln86_87_fu_7628_p2;
wire   [0:0] xor_ln86_64_fu_7640_p2;
wire   [0:0] xor_ln86_63_fu_7634_p2;
wire   [0:0] and_ln87_85_fu_7658_p2;
wire   [0:0] xor_ln87_105_fu_7676_p2;
wire   [0:0] and_ln87_84_fu_7652_p2;
wire   [0:0] and_ln87_87_fu_7670_p2;
wire   [0:0] xor_ln87_107_fu_7688_p2;
wire   [0:0] and_ln87_86_fu_7664_p2;
wire   [0:0] xor_ln87_108_fu_7694_p2;
wire   [0:0] xor_ln87_106_fu_7682_p2;
wire   [0:0] and_ln88_85_fu_7712_p2;
wire   [0:0] and_ln88_86_fu_7718_p2;
wire   [0:0] xor_ln88_105_fu_7730_p2;
wire   [0:0] and_ln88_84_fu_7706_p2;
wire   [0:0] and_ln88_87_fu_7724_p2;
wire   [0:0] xor_ln88_107_fu_7742_p2;
wire   [0:0] xor_ln88_108_fu_7748_p2;
wire   [0:0] xor_ln88_106_fu_7736_p2;
wire   [0:0] and_ln90_63_fu_7760_p2;
wire   [0:0] and_ln90_64_fu_7766_p2;
wire   [0:0] and_ln90_65_fu_7772_p2;
wire   [0:0] xor_ln91_175_fu_7790_p2;
wire   [0:0] xor_ln91_174_fu_7784_p2;
wire   [0:0] xor_ln91_178_fu_7808_p2;
wire   [0:0] and_ln91_21_fu_7778_p2;
wire   [0:0] xor_ln91_179_fu_7814_p2;
wire   [0:0] xor_ln91_177_fu_7802_p2;
wire   [0:0] xor_ln91_180_fu_7820_p2;
wire   [0:0] xor_ln91_176_fu_7796_p2;
wire   [0:0] xor_ln91_43_fu_7826_p2;
wire   [0:0] xor_ln88_109_fu_7754_p2;
wire   [0:0] xor_ln87_109_fu_7700_p2;
wire   [0:0] xor_ln86_65_fu_7646_p2;
wire   [3:0] a0_20_fu_7502_p4;
wire   [3:0] a1_21_fu_7534_p4;
wire   [3:0] xor_ln99_24_fu_7844_p2;
wire   [3:0] b0_9_fu_7518_p4;
wire   [3:0] b1_21_fu_7544_p4;
wire   [3:0] xor_ln99_26_fu_7856_p2;
wire   [3:0] a_40_fu_7850_p2;
wire   [3:0] b_31_fu_7862_p2;
wire   [0:0] trunc_ln86_24_fu_7868_p1;
wire   [0:0] trunc_ln86_25_fu_7872_p1;
wire   [0:0] tmp_164_fu_7882_p3;
wire   [0:0] tmp_165_fu_7890_p3;
wire   [0:0] tmp_166_fu_7904_p3;
wire   [0:0] tmp_167_fu_7912_p3;
wire   [0:0] tmp_168_fu_7926_p3;
wire   [0:0] tmp_169_fu_7934_p3;
wire   [0:0] and_ln86_88_fu_7876_p2;
wire   [0:0] and_ln86_89_fu_7898_p2;
wire   [0:0] and_ln86_90_fu_7920_p2;
wire   [0:0] and_ln86_91_fu_7942_p2;
wire   [0:0] xor_ln86_67_fu_7954_p2;
wire   [0:0] xor_ln86_66_fu_7948_p2;
wire   [0:0] and_ln87_89_fu_7972_p2;
wire   [0:0] xor_ln87_110_fu_7990_p2;
wire   [0:0] and_ln87_88_fu_7966_p2;
wire   [0:0] and_ln87_91_fu_7984_p2;
wire   [0:0] xor_ln87_112_fu_8002_p2;
wire   [0:0] and_ln87_90_fu_7978_p2;
wire   [0:0] xor_ln87_113_fu_8008_p2;
wire   [0:0] xor_ln87_111_fu_7996_p2;
wire   [0:0] and_ln88_89_fu_8026_p2;
wire   [0:0] and_ln88_90_fu_8032_p2;
wire   [0:0] xor_ln88_110_fu_8044_p2;
wire   [0:0] and_ln88_88_fu_8020_p2;
wire   [0:0] and_ln88_91_fu_8038_p2;
wire   [0:0] xor_ln88_112_fu_8056_p2;
wire   [0:0] xor_ln88_113_fu_8062_p2;
wire   [0:0] xor_ln88_111_fu_8050_p2;
wire   [0:0] and_ln90_66_fu_8074_p2;
wire   [0:0] and_ln90_67_fu_8080_p2;
wire   [0:0] and_ln90_68_fu_8086_p2;
wire   [0:0] xor_ln91_182_fu_8104_p2;
wire   [0:0] xor_ln91_181_fu_8098_p2;
wire   [0:0] xor_ln91_185_fu_8122_p2;
wire   [0:0] and_ln91_22_fu_8092_p2;
wire   [0:0] xor_ln91_186_fu_8128_p2;
wire   [0:0] xor_ln91_184_fu_8116_p2;
wire   [0:0] xor_ln91_187_fu_8134_p2;
wire   [0:0] xor_ln91_183_fu_8110_p2;
wire   [0:0] xor_ln91_45_fu_8140_p2;
wire   [0:0] xor_ln88_114_fu_8068_p2;
wire   [0:0] xor_ln87_114_fu_8014_p2;
wire   [0:0] xor_ln86_68_fu_7960_p2;
wire   [0:0] tmp_170_fu_8158_p3;
wire   [0:0] tmp_171_fu_8166_p3;
wire   [0:0] tmp_172_fu_8180_p3;
wire   [0:0] tmp_173_fu_8188_p3;
wire   [0:0] tmp_174_fu_8202_p3;
wire   [0:0] tmp_175_fu_8210_p3;
wire   [0:0] tmp_176_fu_8224_p3;
wire   [0:0] tmp_177_fu_8232_p3;
wire   [0:0] and_ln86_93_fu_8196_p2;
wire   [0:0] and_ln86_94_fu_8218_p2;
wire   [0:0] and_ln86_92_fu_8174_p2;
wire   [0:0] and_ln86_95_fu_8240_p2;
wire   [0:0] xor_ln86_70_fu_8252_p2;
wire   [0:0] xor_ln86_69_fu_8246_p2;
wire   [0:0] and_ln87_93_fu_8270_p2;
wire   [0:0] and_ln87_92_fu_8264_p2;
wire   [0:0] and_ln87_94_fu_8276_p2;
wire   [0:0] xor_ln87_116_fu_8288_p2;
wire   [0:0] xor_ln87_115_fu_8282_p2;
wire   [0:0] and_ln87_95_fu_8300_p2;
wire   [0:0] xor_ln87_118_fu_8306_p2;
wire   [0:0] xor_ln87_117_fu_8294_p2;
wire   [0:0] and_ln88_94_fu_8330_p2;
wire   [0:0] and_ln88_92_fu_8318_p2;
wire   [0:0] and_ln88_95_fu_8336_p2;
wire   [0:0] xor_ln88_116_fu_8348_p2;
wire   [0:0] and_ln88_93_fu_8324_p2;
wire   [0:0] xor_ln88_117_fu_8354_p2;
wire   [0:0] xor_ln88_115_fu_8342_p2;
wire   [0:0] xor_ln88_118_fu_8360_p2;
wire   [0:0] and_ln91_23_fu_8390_p2;
wire   [0:0] xor_ln91_189_fu_8402_p2;
wire   [0:0] xor_ln91_188_fu_8396_p2;
wire   [0:0] and_ln90_70_fu_8378_p2;
wire   [0:0] and_ln90_69_fu_8372_p2;
wire   [0:0] xor_ln91_192_fu_8420_p2;
wire   [0:0] and_ln90_71_fu_8384_p2;
wire   [0:0] xor_ln91_193_fu_8426_p2;
wire   [0:0] xor_ln91_191_fu_8414_p2;
wire   [0:0] xor_ln91_194_fu_8432_p2;
wire   [0:0] xor_ln91_190_fu_8408_p2;
wire   [0:0] xor_ln91_47_fu_8438_p2;
wire   [0:0] xor_ln88_119_fu_8366_p2;
wire   [0:0] xor_ln87_119_fu_8312_p2;
wire   [0:0] xor_ln86_71_fu_8258_p2;
wire   [0:0] xor_ln54_14_fu_8462_p2;
wire   [0:0] xor_ln54_15_fu_8468_p2;
wire   [0:0] xor_ln53_7_fu_8456_p2;
wire   [3:0] res_62_fu_8146_p5;
wire   [3:0] res_61_fu_7832_p5;
wire   [3:0] res_63_fu_8444_p5;
wire   [3:0] res_33_fu_8474_p5;
wire   [3:0] xor_ln101_35_fu_8492_p2;
wire   [3:0] xor_ln101_34_fu_8486_p2;
wire   [3:0] xor_ln101_36_fu_8498_p2;
wire   [3:0] xor_ln101_37_fu_8504_p2;
wire   [0:0] tmp_178_fu_8538_p3;
wire   [0:0] tmp_179_fu_8546_p3;
wire   [0:0] tmp_180_fu_8560_p3;
wire   [0:0] tmp_181_fu_8568_p3;
wire   [0:0] tmp_182_fu_8582_p3;
wire   [0:0] tmp_183_fu_8590_p3;
wire   [0:0] tmp_184_fu_8604_p3;
wire   [0:0] tmp_185_fu_8612_p3;
wire   [0:0] and_ln86_96_fu_8554_p2;
wire   [0:0] and_ln86_97_fu_8576_p2;
wire   [0:0] and_ln86_98_fu_8598_p2;
wire   [0:0] and_ln86_99_fu_8620_p2;
wire   [0:0] xor_ln86_73_fu_8632_p2;
wire   [0:0] xor_ln86_72_fu_8626_p2;
wire   [0:0] and_ln87_97_fu_8650_p2;
wire   [0:0] xor_ln87_120_fu_8668_p2;
wire   [0:0] and_ln87_96_fu_8644_p2;
wire   [0:0] and_ln87_99_fu_8662_p2;
wire   [0:0] xor_ln87_122_fu_8680_p2;
wire   [0:0] and_ln87_98_fu_8656_p2;
wire   [0:0] xor_ln87_123_fu_8686_p2;
wire   [0:0] xor_ln87_121_fu_8674_p2;
wire   [0:0] and_ln88_97_fu_8704_p2;
wire   [0:0] and_ln88_98_fu_8710_p2;
wire   [0:0] xor_ln88_120_fu_8722_p2;
wire   [0:0] and_ln88_96_fu_8698_p2;
wire   [0:0] and_ln88_99_fu_8716_p2;
wire   [0:0] xor_ln88_122_fu_8734_p2;
wire   [0:0] xor_ln88_123_fu_8740_p2;
wire   [0:0] xor_ln88_121_fu_8728_p2;
wire   [0:0] and_ln90_72_fu_8752_p2;
wire   [0:0] and_ln90_73_fu_8758_p2;
wire   [0:0] and_ln90_74_fu_8764_p2;
wire   [0:0] xor_ln91_196_fu_8782_p2;
wire   [0:0] xor_ln91_195_fu_8776_p2;
wire   [0:0] xor_ln91_199_fu_8800_p2;
wire   [0:0] and_ln91_24_fu_8770_p2;
wire   [0:0] xor_ln91_200_fu_8806_p2;
wire   [0:0] xor_ln91_198_fu_8794_p2;
wire   [0:0] xor_ln91_201_fu_8812_p2;
wire   [0:0] xor_ln91_197_fu_8788_p2;
wire   [0:0] xor_ln91_49_fu_8818_p2;
wire   [0:0] xor_ln88_124_fu_8746_p2;
wire   [0:0] xor_ln87_124_fu_8692_p2;
wire   [0:0] xor_ln86_74_fu_8638_p2;
wire   [3:0] a1_22_fu_8518_p4;
wire   [3:0] b1_22_fu_8528_p4;
wire   [3:0] a_45_fu_8836_p2;
wire   [3:0] b_35_fu_8842_p2;
wire   [0:0] trunc_ln86_26_fu_8848_p1;
wire   [0:0] trunc_ln86_27_fu_8852_p1;
wire   [0:0] tmp_186_fu_8862_p3;
wire   [0:0] tmp_187_fu_8870_p3;
wire   [0:0] tmp_188_fu_8884_p3;
wire   [0:0] tmp_189_fu_8892_p3;
wire   [0:0] tmp_190_fu_8906_p3;
wire   [0:0] tmp_191_fu_8914_p3;
wire   [0:0] and_ln86_100_fu_8856_p2;
wire   [0:0] and_ln86_101_fu_8878_p2;
wire   [0:0] and_ln86_102_fu_8900_p2;
wire   [0:0] and_ln86_103_fu_8922_p2;
wire   [0:0] xor_ln86_76_fu_8934_p2;
wire   [0:0] xor_ln86_75_fu_8928_p2;
wire   [0:0] and_ln87_101_fu_8952_p2;
wire   [0:0] xor_ln87_125_fu_8970_p2;
wire   [0:0] and_ln87_100_fu_8946_p2;
wire   [0:0] and_ln87_103_fu_8964_p2;
wire   [0:0] xor_ln87_127_fu_8982_p2;
wire   [0:0] and_ln87_102_fu_8958_p2;
wire   [0:0] xor_ln87_128_fu_8988_p2;
wire   [0:0] xor_ln87_126_fu_8976_p2;
wire   [0:0] and_ln88_101_fu_9006_p2;
wire   [0:0] and_ln88_102_fu_9012_p2;
wire   [0:0] xor_ln88_125_fu_9024_p2;
wire   [0:0] and_ln88_100_fu_9000_p2;
wire   [0:0] and_ln88_103_fu_9018_p2;
wire   [0:0] xor_ln88_127_fu_9036_p2;
wire   [0:0] xor_ln88_128_fu_9042_p2;
wire   [0:0] xor_ln88_126_fu_9030_p2;
wire   [0:0] and_ln90_75_fu_9054_p2;
wire   [0:0] and_ln90_76_fu_9060_p2;
wire   [0:0] and_ln90_77_fu_9066_p2;
wire   [0:0] xor_ln91_203_fu_9084_p2;
wire   [0:0] xor_ln91_202_fu_9078_p2;
wire   [0:0] xor_ln91_206_fu_9102_p2;
wire   [0:0] and_ln91_25_fu_9072_p2;
wire   [0:0] xor_ln91_207_fu_9108_p2;
wire   [0:0] xor_ln91_205_fu_9096_p2;
wire   [0:0] xor_ln91_208_fu_9114_p2;
wire   [0:0] xor_ln91_204_fu_9090_p2;
wire   [0:0] xor_ln91_51_fu_9120_p2;
wire   [0:0] xor_ln88_129_fu_9048_p2;
wire   [0:0] xor_ln87_129_fu_8994_p2;
wire   [0:0] xor_ln86_77_fu_8940_p2;
wire   [0:0] tmp_192_fu_9138_p3;
wire   [0:0] tmp_193_fu_9146_p3;
wire   [0:0] tmp_194_fu_9160_p3;
wire   [0:0] tmp_195_fu_9168_p3;
wire   [0:0] tmp_196_fu_9182_p3;
wire   [0:0] tmp_197_fu_9190_p3;
wire   [0:0] tmp_198_fu_9204_p3;
wire   [0:0] tmp_199_fu_9212_p3;
wire   [0:0] and_ln86_105_fu_9176_p2;
wire   [0:0] and_ln86_106_fu_9198_p2;
wire   [0:0] and_ln86_104_fu_9154_p2;
wire   [0:0] and_ln86_107_fu_9220_p2;
wire   [0:0] xor_ln86_79_fu_9232_p2;
wire   [0:0] xor_ln86_78_fu_9226_p2;
wire   [0:0] and_ln87_105_fu_9250_p2;
wire   [0:0] and_ln87_104_fu_9244_p2;
wire   [0:0] and_ln87_106_fu_9256_p2;
wire   [0:0] xor_ln87_131_fu_9268_p2;
wire   [0:0] xor_ln87_130_fu_9262_p2;
wire   [0:0] and_ln87_107_fu_9280_p2;
wire   [0:0] xor_ln87_133_fu_9286_p2;
wire   [0:0] xor_ln87_132_fu_9274_p2;
wire   [0:0] and_ln88_106_fu_9310_p2;
wire   [0:0] and_ln88_104_fu_9298_p2;
wire   [0:0] and_ln88_107_fu_9316_p2;
wire   [0:0] xor_ln88_131_fu_9328_p2;
wire   [0:0] and_ln88_105_fu_9304_p2;
wire   [0:0] xor_ln88_132_fu_9334_p2;
wire   [0:0] xor_ln88_130_fu_9322_p2;
wire   [0:0] xor_ln88_133_fu_9340_p2;
wire   [0:0] and_ln91_26_fu_9370_p2;
wire   [0:0] xor_ln91_210_fu_9382_p2;
wire   [0:0] xor_ln91_209_fu_9376_p2;
wire   [0:0] and_ln90_79_fu_9358_p2;
wire   [0:0] and_ln90_78_fu_9352_p2;
wire   [0:0] xor_ln91_213_fu_9400_p2;
wire   [0:0] and_ln90_80_fu_9364_p2;
wire   [0:0] xor_ln91_214_fu_9406_p2;
wire   [0:0] xor_ln91_212_fu_9394_p2;
wire   [0:0] xor_ln91_215_fu_9412_p2;
wire   [0:0] xor_ln91_211_fu_9388_p2;
wire   [0:0] xor_ln91_53_fu_9418_p2;
wire   [0:0] xor_ln88_134_fu_9346_p2;
wire   [0:0] xor_ln87_134_fu_9292_p2;
wire   [0:0] xor_ln86_80_fu_9238_p2;
wire   [0:0] xor_ln54_16_fu_9442_p2;
wire   [0:0] xor_ln54_17_fu_9448_p2;
wire   [0:0] xor_ln53_8_fu_9436_p2;
wire   [3:0] res_64_fu_8824_p5;
wire   [3:0] res_66_fu_9424_p5;
wire   [3:0] res_65_fu_9126_p5;
wire   [3:0] res_37_fu_9454_p5;
wire   [3:0] xor_ln101_39_fu_9472_p2;
wire   [3:0] xor_ln101_38_fu_9466_p2;
wire   [3:0] xor_ln101_40_fu_9478_p2;
wire   [0:0] trunc_ln62_2_fu_9492_p1;
wire   [0:0] tmp_200_fu_9496_p3;
wire   [0:0] tmp_201_fu_9510_p3;
wire   [0:0] tmp_202_fu_9518_p3;
wire   [0:0] trunc_ln64_2_fu_9540_p1;
wire   [0:0] xor_ln64_4_fu_9544_p2;
wire   [0:0] tmp_203_fu_9532_p3;
wire   [0:0] tmp_204_fu_9556_p3;
wire   [0:0] tmp_205_fu_9564_p3;
wire   [0:0] xor_ln65_7_fu_9578_p2;
wire   [0:0] xor_ln65_6_fu_9572_p2;
wire   [0:0] xor_ln65_8_fu_9584_p2;
wire   [0:0] xor_ln64_5_fu_9550_p2;
wire   [0:0] xor_ln63_2_fu_9526_p2;
wire   [0:0] xor_ln62_2_fu_9504_p2;
wire   [7:0] z0_10_fu_7494_p3;
wire   [7:0] z2_5_fu_9484_p3;
wire   [7:0] z1_11_fu_8510_p3;
wire   [7:0] res_38_fu_9590_p6;
wire   [7:0] xor_ln101_42_fu_9610_p2;
wire   [7:0] a0_fu_9604_p2;
wire   [7:0] a1_23_fu_9616_p2;
wire   [0:0] trunc_ln62_3_fu_9630_p1;
wire   [0:0] tmp_206_fu_9634_p3;
wire   [0:0] tmp_207_fu_9648_p3;
wire   [0:0] tmp_208_fu_9656_p3;
wire   [0:0] tmp_210_fu_9678_p3;
wire   [0:0] xor_ln64_6_fu_9686_p2;
wire   [0:0] tmp_209_fu_9670_p3;
wire   [0:0] tmp_211_fu_9698_p3;
wire   [0:0] tmp_212_fu_9706_p3;
wire   [0:0] xor_ln65_10_fu_9720_p2;
wire   [0:0] xor_ln65_9_fu_9714_p2;
wire   [0:0] xor_ln65_11_fu_9726_p2;
wire   [0:0] xor_ln64_7_fu_9692_p2;
wire   [0:0] xor_ln63_3_fu_9664_p2;
wire   [0:0] xor_ln62_3_fu_9642_p2;
wire   [3:0] tmp_s_fu_9732_p4;
wire   [7:0] res_39_fu_9742_p6;
wire   [7:0] xor_ln70_fu_9756_p2;
wire   [15:0] z1_8_fu_6494_p3;
wire   [15:0] z0_4_fu_3292_p3;
wire   [15:0] z2_6_fu_9622_p3;
wire   [15:0] tmp_213_fu_9762_p3;
wire   [15:0] xor_ln101_45_fu_9776_p2;
wire   [15:0] xor_ln101_44_fu_9770_p2;
wire   [15:0] xor_ln101_46_fu_9782_p2;
wire   [15:0] xor_ln101_47_fu_9788_p2;

assign a0_11_fu_130_p1 = a[15:0];

assign a0_12_fu_158_p1 = a[7:0];

assign a0_13_fu_186_p1 = a[3:0];

assign a0_14_fu_1166_p4 = {{a[11:8]}};

assign a0_15_fu_3352_p2 = (a0_18_fu_3310_p4 ^ a0_12_fu_158_p1);

assign a0_16_fu_3384_p2 = (a0_19_fu_3300_p4 ^ a0_13_fu_186_p1);

assign a0_17_fu_4368_p4 = {{a_17_fu_3320_p2[11:8]}};

assign a0_18_fu_3310_p4 = {{a[23:16]}};

assign a0_19_fu_3300_p4 = {{a[19:16]}};

assign a0_20_fu_7502_p4 = {{a[27:24]}};

assign a0_fu_9604_p2 = (z2_5_fu_9484_p3 ^ z0_10_fu_7494_p3);

assign a1_11_fu_162_p4 = {{a[15:8]}};

assign a1_12_fu_190_p4 = {{a[7:4]}};

assign a1_13_fu_1198_p4 = {{a_7_fu_1176_p2[7:4]}};

assign a1_14_fu_2182_p4 = {{a[15:12]}};

assign a1_15_fu_3358_p4 = {{a_17_fu_3320_p2[15:8]}};

assign a1_16_fu_3390_p4 = {{a0_15_fu_3352_p2[7:4]}};

assign a1_17_fu_4400_p4 = {{a_23_fu_4378_p2[7:4]}};

assign a1_18_fu_5384_p4 = {{a_17_fu_3320_p2[15:12]}};

assign a1_19_fu_6502_p4 = {{a[31:24]}};

assign a1_20_fu_6522_p4 = {{a[23:20]}};

assign a1_21_fu_7534_p4 = {{a_39_fu_7512_p2[7:4]}};

assign a1_22_fu_8518_p4 = {{a[31:28]}};

assign a1_23_fu_9616_p2 = (xor_ln101_42_fu_9610_p2 ^ a0_fu_9604_p2);

assign a1_fu_134_p4 = {{a[31:16]}};

assign a_13_fu_2500_p2 = (a1_14_fu_2182_p4 ^ a0_14_fu_1166_p4);

assign a_17_fu_3320_p2 = (a1_fu_134_p4 ^ a0_11_fu_130_p1);

assign a_20_fu_3706_p2 = (a1_16_fu_3390_p4 ^ a0_16_fu_3384_p2);

assign a_23_fu_4378_p2 = (a1_15_fu_3358_p4 ^ a0_15_fu_3352_p2);

assign a_24_fu_4716_p2 = (xor_ln99_14_fu_4710_p2 ^ a0_17_fu_4368_p4);

assign a_29_fu_5702_p2 = (a1_18_fu_5384_p4 ^ a0_17_fu_4368_p4);

assign a_36_fu_6840_p2 = (a1_20_fu_6522_p4 ^ a0_19_fu_3300_p4);

assign a_39_fu_7512_p2 = (a1_19_fu_6502_p4 ^ a0_18_fu_3310_p4);

assign a_40_fu_7850_p2 = (xor_ln99_24_fu_7844_p2 ^ a0_19_fu_3300_p4);

assign a_45_fu_8836_p2 = (a1_22_fu_8518_p4 ^ a0_20_fu_7502_p4);

assign a_4_fu_504_p2 = (a1_12_fu_190_p4 ^ a0_13_fu_186_p1);

assign a_7_fu_1176_p2 = (a1_11_fu_162_p4 ^ a0_12_fu_158_p1);

assign a_8_fu_1514_p2 = (xor_ln99_fu_1508_p2 ^ a0_14_fu_1166_p4);

assign and_ln86_100_fu_8856_p2 = (trunc_ln86_27_fu_8852_p1 & trunc_ln86_26_fu_8848_p1);

assign and_ln86_101_fu_8878_p2 = (tmp_187_fu_8870_p3 & tmp_186_fu_8862_p3);

assign and_ln86_102_fu_8900_p2 = (tmp_189_fu_8892_p3 & tmp_188_fu_8884_p3);

assign and_ln86_103_fu_8922_p2 = (tmp_191_fu_8914_p3 & tmp_190_fu_8906_p3);

assign and_ln86_104_fu_9154_p2 = (tmp_193_fu_9146_p3 & tmp_192_fu_9138_p3);

assign and_ln86_105_fu_9176_p2 = (tmp_195_fu_9168_p3 & tmp_194_fu_9160_p3);

assign and_ln86_106_fu_9198_p2 = (tmp_197_fu_9190_p3 & tmp_196_fu_9182_p3);

assign and_ln86_107_fu_9220_p2 = (tmp_199_fu_9212_p3 & tmp_198_fu_9204_p3);

assign and_ln86_10_fu_866_p2 = (tmp_17_fu_858_p3 & tmp_16_fu_850_p3);

assign and_ln86_11_fu_888_p2 = (tmp_19_fu_880_p3 & tmp_18_fu_872_p3);

assign and_ln86_12_fu_1226_p2 = (trunc_ln86_5_fu_1222_p1 & trunc_ln86_4_fu_1218_p1);

assign and_ln86_13_fu_1248_p2 = (tmp_21_fu_1240_p3 & tmp_20_fu_1232_p3);

assign and_ln86_14_fu_1270_p2 = (tmp_23_fu_1262_p3 & tmp_22_fu_1254_p3);

assign and_ln86_15_fu_1292_p2 = (tmp_25_fu_1284_p3 & tmp_24_fu_1276_p3);

assign and_ln86_16_fu_1540_p2 = (trunc_ln86_7_fu_1536_p1 & trunc_ln86_6_fu_1532_p1);

assign and_ln86_17_fu_1562_p2 = (tmp_27_fu_1554_p3 & tmp_26_fu_1546_p3);

assign and_ln86_18_fu_1584_p2 = (tmp_29_fu_1576_p3 & tmp_28_fu_1568_p3);

assign and_ln86_19_fu_1606_p2 = (tmp_31_fu_1598_p3 & tmp_30_fu_1590_p3);

assign and_ln86_1_fu_244_p2 = (tmp_fu_228_p3 & tmp_1_fu_236_p3);

assign and_ln86_20_fu_1838_p2 = (tmp_33_fu_1830_p3 & tmp_32_fu_1822_p3);

assign and_ln86_21_fu_1860_p2 = (tmp_35_fu_1852_p3 & tmp_34_fu_1844_p3);

assign and_ln86_22_fu_1882_p2 = (tmp_37_fu_1874_p3 & tmp_36_fu_1866_p3);

assign and_ln86_23_fu_1904_p2 = (tmp_39_fu_1896_p3 & tmp_38_fu_1888_p3);

assign and_ln86_24_fu_2218_p2 = (tmp_41_fu_2210_p3 & tmp_40_fu_2202_p3);

assign and_ln86_25_fu_2240_p2 = (tmp_43_fu_2232_p3 & tmp_42_fu_2224_p3);

assign and_ln86_26_fu_2262_p2 = (tmp_45_fu_2254_p3 & tmp_44_fu_2246_p3);

assign and_ln86_27_fu_2284_p2 = (tmp_47_fu_2276_p3 & tmp_46_fu_2268_p3);

assign and_ln86_28_fu_2520_p2 = (trunc_ln86_9_fu_2516_p1 & trunc_ln86_8_fu_2512_p1);

assign and_ln86_29_fu_2542_p2 = (tmp_49_fu_2534_p3 & tmp_48_fu_2526_p3);

assign and_ln86_2_fu_266_p2 = (tmp_3_fu_258_p3 & tmp_2_fu_250_p3);

assign and_ln86_30_fu_2564_p2 = (tmp_51_fu_2556_p3 & tmp_50_fu_2548_p3);

assign and_ln86_31_fu_2586_p2 = (tmp_53_fu_2578_p3 & tmp_52_fu_2570_p3);

assign and_ln86_32_fu_2818_p2 = (tmp_55_fu_2810_p3 & tmp_54_fu_2802_p3);

assign and_ln86_33_fu_2840_p2 = (tmp_57_fu_2832_p3 & tmp_56_fu_2824_p3);

assign and_ln86_34_fu_2862_p2 = (tmp_59_fu_2854_p3 & tmp_58_fu_2846_p3);

assign and_ln86_35_fu_2884_p2 = (tmp_61_fu_2876_p3 & tmp_60_fu_2868_p3);

assign and_ln86_36_fu_3424_p2 = (trunc_ln86_11_fu_3420_p1 & trunc_ln86_10_fu_3416_p1);

assign and_ln86_37_fu_3446_p2 = (tmp_69_fu_3438_p3 & tmp_68_fu_3430_p3);

assign and_ln86_38_fu_3468_p2 = (tmp_71_fu_3460_p3 & tmp_70_fu_3452_p3);

assign and_ln86_39_fu_3490_p2 = (tmp_73_fu_3482_p3 & tmp_72_fu_3474_p3);

assign and_ln86_3_fu_288_p2 = (tmp_5_fu_280_p3 & tmp_4_fu_272_p3);

assign and_ln86_40_fu_3726_p2 = (trunc_ln86_13_fu_3722_p1 & trunc_ln86_12_fu_3718_p1);

assign and_ln86_41_fu_3748_p2 = (tmp_75_fu_3740_p3 & tmp_74_fu_3732_p3);

assign and_ln86_42_fu_3770_p2 = (tmp_77_fu_3762_p3 & tmp_76_fu_3754_p3);

assign and_ln86_43_fu_3792_p2 = (tmp_79_fu_3784_p3 & tmp_78_fu_3776_p3);

assign and_ln86_44_fu_4024_p2 = (tmp_81_fu_4016_p3 & tmp_80_fu_4008_p3);

assign and_ln86_45_fu_4046_p2 = (tmp_83_fu_4038_p3 & tmp_82_fu_4030_p3);

assign and_ln86_46_fu_4068_p2 = (tmp_85_fu_4060_p3 & tmp_84_fu_4052_p3);

assign and_ln86_47_fu_4090_p2 = (tmp_87_fu_4082_p3 & tmp_86_fu_4074_p3);

assign and_ln86_48_fu_4428_p2 = (trunc_ln86_15_fu_4424_p1 & trunc_ln86_14_fu_4420_p1);

assign and_ln86_49_fu_4450_p2 = (tmp_89_fu_4442_p3 & tmp_88_fu_4434_p3);

assign and_ln86_4_fu_524_p2 = (trunc_ln86_3_fu_520_p1 & trunc_ln86_2_fu_516_p1);

assign and_ln86_50_fu_4472_p2 = (tmp_91_fu_4464_p3 & tmp_90_fu_4456_p3);

assign and_ln86_51_fu_4494_p2 = (tmp_93_fu_4486_p3 & tmp_92_fu_4478_p3);

assign and_ln86_52_fu_4742_p2 = (trunc_ln86_17_fu_4738_p1 & trunc_ln86_16_fu_4734_p1);

assign and_ln86_53_fu_4764_p2 = (tmp_95_fu_4756_p3 & tmp_94_fu_4748_p3);

assign and_ln86_54_fu_4786_p2 = (tmp_97_fu_4778_p3 & tmp_96_fu_4770_p3);

assign and_ln86_55_fu_4808_p2 = (tmp_99_fu_4800_p3 & tmp_98_fu_4792_p3);

assign and_ln86_56_fu_5040_p2 = (tmp_101_fu_5032_p3 & tmp_100_fu_5024_p3);

assign and_ln86_57_fu_5062_p2 = (tmp_103_fu_5054_p3 & tmp_102_fu_5046_p3);

assign and_ln86_58_fu_5084_p2 = (tmp_105_fu_5076_p3 & tmp_104_fu_5068_p3);

assign and_ln86_59_fu_5106_p2 = (tmp_107_fu_5098_p3 & tmp_106_fu_5090_p3);

assign and_ln86_5_fu_546_p2 = (tmp_7_fu_538_p3 & tmp_6_fu_530_p3);

assign and_ln86_60_fu_5420_p2 = (tmp_109_fu_5412_p3 & tmp_108_fu_5404_p3);

assign and_ln86_61_fu_5442_p2 = (tmp_111_fu_5434_p3 & tmp_110_fu_5426_p3);

assign and_ln86_62_fu_5464_p2 = (tmp_113_fu_5456_p3 & tmp_112_fu_5448_p3);

assign and_ln86_63_fu_5486_p2 = (tmp_115_fu_5478_p3 & tmp_114_fu_5470_p3);

assign and_ln86_64_fu_5722_p2 = (trunc_ln86_19_fu_5718_p1 & trunc_ln86_18_fu_5714_p1);

assign and_ln86_65_fu_5744_p2 = (tmp_117_fu_5736_p3 & tmp_116_fu_5728_p3);

assign and_ln86_66_fu_5766_p2 = (tmp_119_fu_5758_p3 & tmp_118_fu_5750_p3);

assign and_ln86_67_fu_5788_p2 = (tmp_121_fu_5780_p3 & tmp_120_fu_5772_p3);

assign and_ln86_68_fu_6020_p2 = (tmp_123_fu_6012_p3 & tmp_122_fu_6004_p3);

assign and_ln86_69_fu_6042_p2 = (tmp_125_fu_6034_p3 & tmp_124_fu_6026_p3);

assign and_ln86_6_fu_568_p2 = (tmp_9_fu_560_p3 & tmp_8_fu_552_p3);

assign and_ln86_70_fu_6064_p2 = (tmp_127_fu_6056_p3 & tmp_126_fu_6048_p3);

assign and_ln86_71_fu_6086_p2 = (tmp_129_fu_6078_p3 & tmp_128_fu_6070_p3);

assign and_ln86_72_fu_6558_p2 = (tmp_137_fu_6550_p3 & tmp_136_fu_6542_p3);

assign and_ln86_73_fu_6580_p2 = (tmp_139_fu_6572_p3 & tmp_138_fu_6564_p3);

assign and_ln86_74_fu_6602_p2 = (tmp_141_fu_6594_p3 & tmp_140_fu_6586_p3);

assign and_ln86_75_fu_6624_p2 = (tmp_143_fu_6616_p3 & tmp_142_fu_6608_p3);

assign and_ln86_76_fu_6860_p2 = (trunc_ln86_21_fu_6856_p1 & trunc_ln86_20_fu_6852_p1);

assign and_ln86_77_fu_6882_p2 = (tmp_145_fu_6874_p3 & tmp_144_fu_6866_p3);

assign and_ln86_78_fu_6904_p2 = (tmp_147_fu_6896_p3 & tmp_146_fu_6888_p3);

assign and_ln86_79_fu_6926_p2 = (tmp_149_fu_6918_p3 & tmp_148_fu_6910_p3);

assign and_ln86_7_fu_590_p2 = (tmp_11_fu_582_p3 & tmp_10_fu_574_p3);

assign and_ln86_80_fu_7158_p2 = (tmp_151_fu_7150_p3 & tmp_150_fu_7142_p3);

assign and_ln86_81_fu_7180_p2 = (tmp_153_fu_7172_p3 & tmp_152_fu_7164_p3);

assign and_ln86_82_fu_7202_p2 = (tmp_155_fu_7194_p3 & tmp_154_fu_7186_p3);

assign and_ln86_83_fu_7224_p2 = (tmp_157_fu_7216_p3 & tmp_156_fu_7208_p3);

assign and_ln86_84_fu_7562_p2 = (trunc_ln86_23_fu_7558_p1 & trunc_ln86_22_fu_7554_p1);

assign and_ln86_85_fu_7584_p2 = (tmp_159_fu_7576_p3 & tmp_158_fu_7568_p3);

assign and_ln86_86_fu_7606_p2 = (tmp_161_fu_7598_p3 & tmp_160_fu_7590_p3);

assign and_ln86_87_fu_7628_p2 = (tmp_163_fu_7620_p3 & tmp_162_fu_7612_p3);

assign and_ln86_88_fu_7876_p2 = (trunc_ln86_25_fu_7872_p1 & trunc_ln86_24_fu_7868_p1);

assign and_ln86_89_fu_7898_p2 = (tmp_165_fu_7890_p3 & tmp_164_fu_7882_p3);

assign and_ln86_8_fu_822_p2 = (tmp_13_fu_814_p3 & tmp_12_fu_806_p3);

assign and_ln86_90_fu_7920_p2 = (tmp_167_fu_7912_p3 & tmp_166_fu_7904_p3);

assign and_ln86_91_fu_7942_p2 = (tmp_169_fu_7934_p3 & tmp_168_fu_7926_p3);

assign and_ln86_92_fu_8174_p2 = (tmp_171_fu_8166_p3 & tmp_170_fu_8158_p3);

assign and_ln86_93_fu_8196_p2 = (tmp_173_fu_8188_p3 & tmp_172_fu_8180_p3);

assign and_ln86_94_fu_8218_p2 = (tmp_175_fu_8210_p3 & tmp_174_fu_8202_p3);

assign and_ln86_95_fu_8240_p2 = (tmp_177_fu_8232_p3 & tmp_176_fu_8224_p3);

assign and_ln86_96_fu_8554_p2 = (tmp_179_fu_8546_p3 & tmp_178_fu_8538_p3);

assign and_ln86_97_fu_8576_p2 = (tmp_181_fu_8568_p3 & tmp_180_fu_8560_p3);

assign and_ln86_98_fu_8598_p2 = (tmp_183_fu_8590_p3 & tmp_182_fu_8582_p3);

assign and_ln86_99_fu_8620_p2 = (tmp_185_fu_8612_p3 & tmp_184_fu_8604_p3);

assign and_ln86_9_fu_844_p2 = (tmp_15_fu_836_p3 & tmp_14_fu_828_p3);

assign and_ln86_fu_222_p2 = (trunc_ln86_fu_214_p1 & trunc_ln86_1_fu_218_p1);

assign and_ln87_100_fu_8946_p2 = (trunc_ln86_27_fu_8852_p1 & tmp_186_fu_8862_p3);

assign and_ln87_101_fu_8952_p2 = (trunc_ln86_26_fu_8848_p1 & tmp_187_fu_8870_p3);

assign and_ln87_102_fu_8958_p2 = (tmp_190_fu_8906_p3 & tmp_189_fu_8892_p3);

assign and_ln87_103_fu_8964_p2 = (tmp_191_fu_8914_p3 & tmp_188_fu_8884_p3);

assign and_ln87_104_fu_9244_p2 = (tmp_194_fu_9160_p3 & tmp_193_fu_9146_p3);

assign and_ln87_105_fu_9250_p2 = (tmp_195_fu_9168_p3 & tmp_192_fu_9138_p3);

assign and_ln87_106_fu_9256_p2 = (tmp_198_fu_9204_p3 & tmp_197_fu_9190_p3);

assign and_ln87_107_fu_9280_p2 = (tmp_199_fu_9212_p3 & tmp_196_fu_9182_p3);

assign and_ln87_10_fu_924_p2 = (tmp_18_fu_872_p3 & tmp_17_fu_858_p3);

assign and_ln87_11_fu_948_p2 = (tmp_19_fu_880_p3 & tmp_16_fu_850_p3);

assign and_ln87_12_fu_1316_p2 = (trunc_ln86_5_fu_1222_p1 & tmp_20_fu_1232_p3);

assign and_ln87_13_fu_1322_p2 = (trunc_ln86_4_fu_1218_p1 & tmp_21_fu_1240_p3);

assign and_ln87_14_fu_1328_p2 = (tmp_24_fu_1276_p3 & tmp_23_fu_1262_p3);

assign and_ln87_15_fu_1334_p2 = (tmp_25_fu_1284_p3 & tmp_22_fu_1254_p3);

assign and_ln87_16_fu_1630_p2 = (trunc_ln86_7_fu_1536_p1 & tmp_26_fu_1546_p3);

assign and_ln87_17_fu_1636_p2 = (trunc_ln86_6_fu_1532_p1 & tmp_27_fu_1554_p3);

assign and_ln87_18_fu_1642_p2 = (tmp_30_fu_1590_p3 & tmp_29_fu_1576_p3);

assign and_ln87_19_fu_1648_p2 = (tmp_31_fu_1598_p3 & tmp_28_fu_1568_p3);

assign and_ln87_1_fu_318_p2 = (trunc_ln86_fu_214_p1 & tmp_1_fu_236_p3);

assign and_ln87_20_fu_1928_p2 = (tmp_34_fu_1844_p3 & tmp_33_fu_1830_p3);

assign and_ln87_21_fu_1934_p2 = (tmp_35_fu_1852_p3 & tmp_32_fu_1822_p3);

assign and_ln87_22_fu_1940_p2 = (tmp_38_fu_1888_p3 & tmp_37_fu_1874_p3);

assign and_ln87_23_fu_1964_p2 = (tmp_39_fu_1896_p3 & tmp_36_fu_1866_p3);

assign and_ln87_24_fu_2308_p2 = (tmp_42_fu_2224_p3 & tmp_41_fu_2210_p3);

assign and_ln87_25_fu_2314_p2 = (tmp_43_fu_2232_p3 & tmp_40_fu_2202_p3);

assign and_ln87_26_fu_2320_p2 = (tmp_46_fu_2268_p3 & tmp_45_fu_2254_p3);

assign and_ln87_27_fu_2326_p2 = (tmp_47_fu_2276_p3 & tmp_44_fu_2246_p3);

assign and_ln87_28_fu_2610_p2 = (trunc_ln86_9_fu_2516_p1 & tmp_48_fu_2526_p3);

assign and_ln87_29_fu_2616_p2 = (trunc_ln86_8_fu_2512_p1 & tmp_49_fu_2534_p3);

assign and_ln87_2_fu_324_p2 = (tmp_4_fu_272_p3 & tmp_3_fu_258_p3);

assign and_ln87_30_fu_2622_p2 = (tmp_52_fu_2570_p3 & tmp_51_fu_2556_p3);

assign and_ln87_31_fu_2628_p2 = (tmp_53_fu_2578_p3 & tmp_50_fu_2548_p3);

assign and_ln87_32_fu_2908_p2 = (tmp_56_fu_2824_p3 & tmp_55_fu_2810_p3);

assign and_ln87_33_fu_2914_p2 = (tmp_57_fu_2832_p3 & tmp_54_fu_2802_p3);

assign and_ln87_34_fu_2920_p2 = (tmp_60_fu_2868_p3 & tmp_59_fu_2854_p3);

assign and_ln87_35_fu_2944_p2 = (tmp_61_fu_2876_p3 & tmp_58_fu_2846_p3);

assign and_ln87_36_fu_3514_p2 = (trunc_ln86_11_fu_3420_p1 & tmp_68_fu_3430_p3);

assign and_ln87_37_fu_3520_p2 = (trunc_ln86_10_fu_3416_p1 & tmp_69_fu_3438_p3);

assign and_ln87_38_fu_3526_p2 = (tmp_72_fu_3474_p3 & tmp_71_fu_3460_p3);

assign and_ln87_39_fu_3532_p2 = (tmp_73_fu_3482_p3 & tmp_70_fu_3452_p3);

assign and_ln87_3_fu_330_p2 = (tmp_5_fu_280_p3 & tmp_2_fu_250_p3);

assign and_ln87_40_fu_3816_p2 = (trunc_ln86_13_fu_3722_p1 & tmp_74_fu_3732_p3);

assign and_ln87_41_fu_3822_p2 = (trunc_ln86_12_fu_3718_p1 & tmp_75_fu_3740_p3);

assign and_ln87_42_fu_3828_p2 = (tmp_78_fu_3776_p3 & tmp_77_fu_3762_p3);

assign and_ln87_43_fu_3834_p2 = (tmp_79_fu_3784_p3 & tmp_76_fu_3754_p3);

assign and_ln87_44_fu_4114_p2 = (tmp_82_fu_4030_p3 & tmp_81_fu_4016_p3);

assign and_ln87_45_fu_4120_p2 = (tmp_83_fu_4038_p3 & tmp_80_fu_4008_p3);

assign and_ln87_46_fu_4126_p2 = (tmp_86_fu_4074_p3 & tmp_85_fu_4060_p3);

assign and_ln87_47_fu_4150_p2 = (tmp_87_fu_4082_p3 & tmp_84_fu_4052_p3);

assign and_ln87_48_fu_4518_p2 = (trunc_ln86_15_fu_4424_p1 & tmp_88_fu_4434_p3);

assign and_ln87_49_fu_4524_p2 = (trunc_ln86_14_fu_4420_p1 & tmp_89_fu_4442_p3);

assign and_ln87_4_fu_614_p2 = (trunc_ln86_3_fu_520_p1 & tmp_6_fu_530_p3);

assign and_ln87_50_fu_4530_p2 = (tmp_92_fu_4478_p3 & tmp_91_fu_4464_p3);

assign and_ln87_51_fu_4536_p2 = (tmp_93_fu_4486_p3 & tmp_90_fu_4456_p3);

assign and_ln87_52_fu_4832_p2 = (trunc_ln86_17_fu_4738_p1 & tmp_94_fu_4748_p3);

assign and_ln87_53_fu_4838_p2 = (trunc_ln86_16_fu_4734_p1 & tmp_95_fu_4756_p3);

assign and_ln87_54_fu_4844_p2 = (tmp_98_fu_4792_p3 & tmp_97_fu_4778_p3);

assign and_ln87_55_fu_4850_p2 = (tmp_99_fu_4800_p3 & tmp_96_fu_4770_p3);

assign and_ln87_56_fu_5130_p2 = (tmp_102_fu_5046_p3 & tmp_101_fu_5032_p3);

assign and_ln87_57_fu_5136_p2 = (tmp_103_fu_5054_p3 & tmp_100_fu_5024_p3);

assign and_ln87_58_fu_5142_p2 = (tmp_106_fu_5090_p3 & tmp_105_fu_5076_p3);

assign and_ln87_59_fu_5166_p2 = (tmp_107_fu_5098_p3 & tmp_104_fu_5068_p3);

assign and_ln87_5_fu_620_p2 = (trunc_ln86_2_fu_516_p1 & tmp_7_fu_538_p3);

assign and_ln87_60_fu_5510_p2 = (tmp_110_fu_5426_p3 & tmp_109_fu_5412_p3);

assign and_ln87_61_fu_5516_p2 = (tmp_111_fu_5434_p3 & tmp_108_fu_5404_p3);

assign and_ln87_62_fu_5522_p2 = (tmp_114_fu_5470_p3 & tmp_113_fu_5456_p3);

assign and_ln87_63_fu_5528_p2 = (tmp_115_fu_5478_p3 & tmp_112_fu_5448_p3);

assign and_ln87_64_fu_5812_p2 = (trunc_ln86_19_fu_5718_p1 & tmp_116_fu_5728_p3);

assign and_ln87_65_fu_5818_p2 = (trunc_ln86_18_fu_5714_p1 & tmp_117_fu_5736_p3);

assign and_ln87_66_fu_5824_p2 = (tmp_120_fu_5772_p3 & tmp_119_fu_5758_p3);

assign and_ln87_67_fu_5830_p2 = (tmp_121_fu_5780_p3 & tmp_118_fu_5750_p3);

assign and_ln87_68_fu_6110_p2 = (tmp_124_fu_6026_p3 & tmp_123_fu_6012_p3);

assign and_ln87_69_fu_6116_p2 = (tmp_125_fu_6034_p3 & tmp_122_fu_6004_p3);

assign and_ln87_6_fu_626_p2 = (tmp_9_fu_560_p3 & tmp_10_fu_574_p3);

assign and_ln87_70_fu_6122_p2 = (tmp_128_fu_6070_p3 & tmp_127_fu_6056_p3);

assign and_ln87_71_fu_6146_p2 = (tmp_129_fu_6078_p3 & tmp_126_fu_6048_p3);

assign and_ln87_72_fu_6648_p2 = (tmp_138_fu_6564_p3 & tmp_137_fu_6550_p3);

assign and_ln87_73_fu_6654_p2 = (tmp_139_fu_6572_p3 & tmp_136_fu_6542_p3);

assign and_ln87_74_fu_6660_p2 = (tmp_142_fu_6608_p3 & tmp_141_fu_6594_p3);

assign and_ln87_75_fu_6666_p2 = (tmp_143_fu_6616_p3 & tmp_140_fu_6586_p3);

assign and_ln87_76_fu_6950_p2 = (trunc_ln86_21_fu_6856_p1 & tmp_144_fu_6866_p3);

assign and_ln87_77_fu_6956_p2 = (trunc_ln86_20_fu_6852_p1 & tmp_145_fu_6874_p3);

assign and_ln87_78_fu_6962_p2 = (tmp_148_fu_6910_p3 & tmp_147_fu_6896_p3);

assign and_ln87_79_fu_6968_p2 = (tmp_149_fu_6918_p3 & tmp_146_fu_6888_p3);

assign and_ln87_7_fu_632_p2 = (tmp_8_fu_552_p3 & tmp_11_fu_582_p3);

assign and_ln87_80_fu_7248_p2 = (tmp_152_fu_7164_p3 & tmp_151_fu_7150_p3);

assign and_ln87_81_fu_7254_p2 = (tmp_153_fu_7172_p3 & tmp_150_fu_7142_p3);

assign and_ln87_82_fu_7260_p2 = (tmp_156_fu_7208_p3 & tmp_155_fu_7194_p3);

assign and_ln87_83_fu_7284_p2 = (tmp_157_fu_7216_p3 & tmp_154_fu_7186_p3);

assign and_ln87_84_fu_7652_p2 = (trunc_ln86_23_fu_7558_p1 & tmp_158_fu_7568_p3);

assign and_ln87_85_fu_7658_p2 = (trunc_ln86_22_fu_7554_p1 & tmp_159_fu_7576_p3);

assign and_ln87_86_fu_7664_p2 = (tmp_162_fu_7612_p3 & tmp_161_fu_7598_p3);

assign and_ln87_87_fu_7670_p2 = (tmp_163_fu_7620_p3 & tmp_160_fu_7590_p3);

assign and_ln87_88_fu_7966_p2 = (trunc_ln86_25_fu_7872_p1 & tmp_164_fu_7882_p3);

assign and_ln87_89_fu_7972_p2 = (trunc_ln86_24_fu_7868_p1 & tmp_165_fu_7890_p3);

assign and_ln87_8_fu_912_p2 = (tmp_14_fu_828_p3 & tmp_13_fu_814_p3);

assign and_ln87_90_fu_7978_p2 = (tmp_168_fu_7926_p3 & tmp_167_fu_7912_p3);

assign and_ln87_91_fu_7984_p2 = (tmp_169_fu_7934_p3 & tmp_166_fu_7904_p3);

assign and_ln87_92_fu_8264_p2 = (tmp_172_fu_8180_p3 & tmp_171_fu_8166_p3);

assign and_ln87_93_fu_8270_p2 = (tmp_173_fu_8188_p3 & tmp_170_fu_8158_p3);

assign and_ln87_94_fu_8276_p2 = (tmp_176_fu_8224_p3 & tmp_175_fu_8210_p3);

assign and_ln87_95_fu_8300_p2 = (tmp_177_fu_8232_p3 & tmp_174_fu_8202_p3);

assign and_ln87_96_fu_8644_p2 = (tmp_180_fu_8560_p3 & tmp_179_fu_8546_p3);

assign and_ln87_97_fu_8650_p2 = (tmp_181_fu_8568_p3 & tmp_178_fu_8538_p3);

assign and_ln87_98_fu_8656_p2 = (tmp_184_fu_8604_p3 & tmp_183_fu_8590_p3);

assign and_ln87_99_fu_8662_p2 = (tmp_185_fu_8612_p3 & tmp_182_fu_8582_p3);

assign and_ln87_9_fu_918_p2 = (tmp_15_fu_836_p3 & tmp_12_fu_806_p3);

assign and_ln87_fu_312_p2 = (trunc_ln86_1_fu_218_p1 & tmp_fu_228_p3);

assign and_ln88_100_fu_9000_p2 = (trunc_ln86_27_fu_8852_p1 & tmp_188_fu_8884_p3);

assign and_ln88_101_fu_9006_p2 = (tmp_190_fu_8906_p3 & tmp_187_fu_8870_p3);

assign and_ln88_102_fu_9012_p2 = (trunc_ln86_26_fu_8848_p1 & tmp_189_fu_8892_p3);

assign and_ln88_103_fu_9018_p2 = (tmp_191_fu_8914_p3 & tmp_186_fu_8862_p3);

assign and_ln88_104_fu_9298_p2 = (tmp_196_fu_9182_p3 & tmp_193_fu_9146_p3);

assign and_ln88_105_fu_9304_p2 = (tmp_198_fu_9204_p3 & tmp_195_fu_9168_p3);

assign and_ln88_106_fu_9310_p2 = (tmp_197_fu_9190_p3 & tmp_192_fu_9138_p3);

assign and_ln88_107_fu_9316_p2 = (tmp_199_fu_9212_p3 & tmp_194_fu_9160_p3);

assign and_ln88_10_fu_978_p2 = (tmp_17_fu_858_p3 & tmp_12_fu_806_p3);

assign and_ln88_11_fu_984_p2 = (tmp_19_fu_880_p3 & tmp_14_fu_828_p3);

assign and_ln88_12_fu_1370_p2 = (trunc_ln86_5_fu_1222_p1 & tmp_22_fu_1254_p3);

assign and_ln88_13_fu_1376_p2 = (tmp_24_fu_1276_p3 & tmp_21_fu_1240_p3);

assign and_ln88_14_fu_1382_p2 = (trunc_ln86_4_fu_1218_p1 & tmp_23_fu_1262_p3);

assign and_ln88_15_fu_1388_p2 = (tmp_25_fu_1284_p3 & tmp_20_fu_1232_p3);

assign and_ln88_16_fu_1684_p2 = (trunc_ln86_7_fu_1536_p1 & tmp_28_fu_1568_p3);

assign and_ln88_17_fu_1690_p2 = (tmp_30_fu_1590_p3 & tmp_27_fu_1554_p3);

assign and_ln88_18_fu_1696_p2 = (trunc_ln86_6_fu_1532_p1 & tmp_29_fu_1576_p3);

assign and_ln88_19_fu_1702_p2 = (tmp_31_fu_1598_p3 & tmp_26_fu_1546_p3);

assign and_ln88_1_fu_372_p2 = (tmp_4_fu_272_p3 & tmp_1_fu_236_p3);

assign and_ln88_20_fu_1982_p2 = (tmp_36_fu_1866_p3 & tmp_33_fu_1830_p3);

assign and_ln88_21_fu_1988_p2 = (tmp_38_fu_1888_p3 & tmp_35_fu_1852_p3);

assign and_ln88_22_fu_1994_p2 = (tmp_37_fu_1874_p3 & tmp_32_fu_1822_p3);

assign and_ln88_23_fu_2000_p2 = (tmp_39_fu_1896_p3 & tmp_34_fu_1844_p3);

assign and_ln88_24_fu_2362_p2 = (tmp_44_fu_2246_p3 & tmp_41_fu_2210_p3);

assign and_ln88_25_fu_2368_p2 = (tmp_46_fu_2268_p3 & tmp_43_fu_2232_p3);

assign and_ln88_26_fu_2374_p2 = (tmp_45_fu_2254_p3 & tmp_40_fu_2202_p3);

assign and_ln88_27_fu_2380_p2 = (tmp_47_fu_2276_p3 & tmp_42_fu_2224_p3);

assign and_ln88_28_fu_2664_p2 = (trunc_ln86_9_fu_2516_p1 & tmp_50_fu_2548_p3);

assign and_ln88_29_fu_2670_p2 = (tmp_52_fu_2570_p3 & tmp_49_fu_2534_p3);

assign and_ln88_2_fu_378_p2 = (trunc_ln86_fu_214_p1 & tmp_3_fu_258_p3);

assign and_ln88_30_fu_2676_p2 = (trunc_ln86_8_fu_2512_p1 & tmp_51_fu_2556_p3);

assign and_ln88_31_fu_2682_p2 = (tmp_53_fu_2578_p3 & tmp_48_fu_2526_p3);

assign and_ln88_32_fu_2962_p2 = (tmp_58_fu_2846_p3 & tmp_55_fu_2810_p3);

assign and_ln88_33_fu_2968_p2 = (tmp_60_fu_2868_p3 & tmp_57_fu_2832_p3);

assign and_ln88_34_fu_2974_p2 = (tmp_59_fu_2854_p3 & tmp_54_fu_2802_p3);

assign and_ln88_35_fu_2980_p2 = (tmp_61_fu_2876_p3 & tmp_56_fu_2824_p3);

assign and_ln88_36_fu_3568_p2 = (trunc_ln86_11_fu_3420_p1 & tmp_70_fu_3452_p3);

assign and_ln88_37_fu_3574_p2 = (tmp_72_fu_3474_p3 & tmp_69_fu_3438_p3);

assign and_ln88_38_fu_3580_p2 = (trunc_ln86_10_fu_3416_p1 & tmp_71_fu_3460_p3);

assign and_ln88_39_fu_3586_p2 = (tmp_73_fu_3482_p3 & tmp_68_fu_3430_p3);

assign and_ln88_3_fu_384_p2 = (tmp_fu_228_p3 & tmp_5_fu_280_p3);

assign and_ln88_40_fu_3870_p2 = (trunc_ln86_13_fu_3722_p1 & tmp_76_fu_3754_p3);

assign and_ln88_41_fu_3876_p2 = (tmp_78_fu_3776_p3 & tmp_75_fu_3740_p3);

assign and_ln88_42_fu_3882_p2 = (trunc_ln86_12_fu_3718_p1 & tmp_77_fu_3762_p3);

assign and_ln88_43_fu_3888_p2 = (tmp_79_fu_3784_p3 & tmp_74_fu_3732_p3);

assign and_ln88_44_fu_4168_p2 = (tmp_84_fu_4052_p3 & tmp_81_fu_4016_p3);

assign and_ln88_45_fu_4174_p2 = (tmp_86_fu_4074_p3 & tmp_83_fu_4038_p3);

assign and_ln88_46_fu_4180_p2 = (tmp_85_fu_4060_p3 & tmp_80_fu_4008_p3);

assign and_ln88_47_fu_4186_p2 = (tmp_87_fu_4082_p3 & tmp_82_fu_4030_p3);

assign and_ln88_48_fu_4572_p2 = (trunc_ln86_15_fu_4424_p1 & tmp_90_fu_4456_p3);

assign and_ln88_49_fu_4578_p2 = (tmp_92_fu_4478_p3 & tmp_89_fu_4442_p3);

assign and_ln88_4_fu_668_p2 = (trunc_ln86_3_fu_520_p1 & tmp_8_fu_552_p3);

assign and_ln88_50_fu_4584_p2 = (trunc_ln86_14_fu_4420_p1 & tmp_91_fu_4464_p3);

assign and_ln88_51_fu_4590_p2 = (tmp_93_fu_4486_p3 & tmp_88_fu_4434_p3);

assign and_ln88_52_fu_4886_p2 = (trunc_ln86_17_fu_4738_p1 & tmp_96_fu_4770_p3);

assign and_ln88_53_fu_4892_p2 = (tmp_98_fu_4792_p3 & tmp_95_fu_4756_p3);

assign and_ln88_54_fu_4898_p2 = (trunc_ln86_16_fu_4734_p1 & tmp_97_fu_4778_p3);

assign and_ln88_55_fu_4904_p2 = (tmp_99_fu_4800_p3 & tmp_94_fu_4748_p3);

assign and_ln88_56_fu_5184_p2 = (tmp_104_fu_5068_p3 & tmp_101_fu_5032_p3);

assign and_ln88_57_fu_5190_p2 = (tmp_106_fu_5090_p3 & tmp_103_fu_5054_p3);

assign and_ln88_58_fu_5196_p2 = (tmp_105_fu_5076_p3 & tmp_100_fu_5024_p3);

assign and_ln88_59_fu_5202_p2 = (tmp_107_fu_5098_p3 & tmp_102_fu_5046_p3);

assign and_ln88_5_fu_674_p2 = (tmp_7_fu_538_p3 & tmp_10_fu_574_p3);

assign and_ln88_60_fu_5564_p2 = (tmp_112_fu_5448_p3 & tmp_109_fu_5412_p3);

assign and_ln88_61_fu_5570_p2 = (tmp_114_fu_5470_p3 & tmp_111_fu_5434_p3);

assign and_ln88_62_fu_5576_p2 = (tmp_113_fu_5456_p3 & tmp_108_fu_5404_p3);

assign and_ln88_63_fu_5582_p2 = (tmp_115_fu_5478_p3 & tmp_110_fu_5426_p3);

assign and_ln88_64_fu_5866_p2 = (trunc_ln86_19_fu_5718_p1 & tmp_118_fu_5750_p3);

assign and_ln88_65_fu_5872_p2 = (tmp_120_fu_5772_p3 & tmp_117_fu_5736_p3);

assign and_ln88_66_fu_5878_p2 = (trunc_ln86_18_fu_5714_p1 & tmp_119_fu_5758_p3);

assign and_ln88_67_fu_5884_p2 = (tmp_121_fu_5780_p3 & tmp_116_fu_5728_p3);

assign and_ln88_68_fu_6164_p2 = (tmp_126_fu_6048_p3 & tmp_123_fu_6012_p3);

assign and_ln88_69_fu_6170_p2 = (tmp_128_fu_6070_p3 & tmp_125_fu_6034_p3);

assign and_ln88_6_fu_680_p2 = (trunc_ln86_2_fu_516_p1 & tmp_9_fu_560_p3);

assign and_ln88_70_fu_6176_p2 = (tmp_127_fu_6056_p3 & tmp_122_fu_6004_p3);

assign and_ln88_71_fu_6182_p2 = (tmp_129_fu_6078_p3 & tmp_124_fu_6026_p3);

assign and_ln88_72_fu_6702_p2 = (tmp_140_fu_6586_p3 & tmp_137_fu_6550_p3);

assign and_ln88_73_fu_6708_p2 = (tmp_142_fu_6608_p3 & tmp_139_fu_6572_p3);

assign and_ln88_74_fu_6714_p2 = (tmp_141_fu_6594_p3 & tmp_136_fu_6542_p3);

assign and_ln88_75_fu_6720_p2 = (tmp_143_fu_6616_p3 & tmp_138_fu_6564_p3);

assign and_ln88_76_fu_7004_p2 = (trunc_ln86_21_fu_6856_p1 & tmp_146_fu_6888_p3);

assign and_ln88_77_fu_7010_p2 = (tmp_148_fu_6910_p3 & tmp_145_fu_6874_p3);

assign and_ln88_78_fu_7016_p2 = (trunc_ln86_20_fu_6852_p1 & tmp_147_fu_6896_p3);

assign and_ln88_79_fu_7022_p2 = (tmp_149_fu_6918_p3 & tmp_144_fu_6866_p3);

assign and_ln88_7_fu_686_p2 = (tmp_6_fu_530_p3 & tmp_11_fu_582_p3);

assign and_ln88_80_fu_7302_p2 = (tmp_154_fu_7186_p3 & tmp_151_fu_7150_p3);

assign and_ln88_81_fu_7308_p2 = (tmp_156_fu_7208_p3 & tmp_153_fu_7172_p3);

assign and_ln88_82_fu_7314_p2 = (tmp_155_fu_7194_p3 & tmp_150_fu_7142_p3);

assign and_ln88_83_fu_7320_p2 = (tmp_157_fu_7216_p3 & tmp_152_fu_7164_p3);

assign and_ln88_84_fu_7706_p2 = (trunc_ln86_23_fu_7558_p1 & tmp_160_fu_7590_p3);

assign and_ln88_85_fu_7712_p2 = (tmp_162_fu_7612_p3 & tmp_159_fu_7576_p3);

assign and_ln88_86_fu_7718_p2 = (trunc_ln86_22_fu_7554_p1 & tmp_161_fu_7598_p3);

assign and_ln88_87_fu_7724_p2 = (tmp_163_fu_7620_p3 & tmp_158_fu_7568_p3);

assign and_ln88_88_fu_8020_p2 = (trunc_ln86_25_fu_7872_p1 & tmp_166_fu_7904_p3);

assign and_ln88_89_fu_8026_p2 = (tmp_168_fu_7926_p3 & tmp_165_fu_7890_p3);

assign and_ln88_8_fu_966_p2 = (tmp_16_fu_850_p3 & tmp_13_fu_814_p3);

assign and_ln88_90_fu_8032_p2 = (trunc_ln86_24_fu_7868_p1 & tmp_167_fu_7912_p3);

assign and_ln88_91_fu_8038_p2 = (tmp_169_fu_7934_p3 & tmp_164_fu_7882_p3);

assign and_ln88_92_fu_8318_p2 = (tmp_174_fu_8202_p3 & tmp_171_fu_8166_p3);

assign and_ln88_93_fu_8324_p2 = (tmp_176_fu_8224_p3 & tmp_173_fu_8188_p3);

assign and_ln88_94_fu_8330_p2 = (tmp_175_fu_8210_p3 & tmp_170_fu_8158_p3);

assign and_ln88_95_fu_8336_p2 = (tmp_177_fu_8232_p3 & tmp_172_fu_8180_p3);

assign and_ln88_96_fu_8698_p2 = (tmp_182_fu_8582_p3 & tmp_179_fu_8546_p3);

assign and_ln88_97_fu_8704_p2 = (tmp_184_fu_8604_p3 & tmp_181_fu_8568_p3);

assign and_ln88_98_fu_8710_p2 = (tmp_183_fu_8590_p3 & tmp_178_fu_8538_p3);

assign and_ln88_99_fu_8716_p2 = (tmp_185_fu_8612_p3 & tmp_180_fu_8560_p3);

assign and_ln88_9_fu_972_p2 = (tmp_18_fu_872_p3 & tmp_15_fu_836_p3);

assign and_ln88_fu_366_p2 = (trunc_ln86_1_fu_218_p1 & tmp_2_fu_250_p3);

assign and_ln90_10_fu_1430_p2 = (tmp_22_fu_1254_p3 & tmp_21_fu_1240_p3);

assign and_ln90_11_fu_1436_p2 = (tmp_23_fu_1262_p3 & tmp_20_fu_1232_p3);

assign and_ln90_12_fu_1738_p2 = (trunc_ln86_7_fu_1536_p1 & tmp_30_fu_1590_p3);

assign and_ln90_13_fu_1744_p2 = (tmp_28_fu_1568_p3 & tmp_27_fu_1554_p3);

assign and_ln90_14_fu_1750_p2 = (tmp_29_fu_1576_p3 & tmp_26_fu_1546_p3);

assign and_ln90_15_fu_2036_p2 = (tmp_38_fu_1888_p3 & tmp_33_fu_1830_p3);

assign and_ln90_16_fu_2042_p2 = (tmp_36_fu_1866_p3 & tmp_35_fu_1852_p3);

assign and_ln90_17_fu_2048_p2 = (tmp_37_fu_1874_p3 & tmp_34_fu_1844_p3);

assign and_ln90_18_fu_2416_p2 = (tmp_46_fu_2268_p3 & tmp_41_fu_2210_p3);

assign and_ln90_19_fu_2422_p2 = (tmp_44_fu_2246_p3 & tmp_43_fu_2232_p3);

assign and_ln90_1_fu_426_p2 = (tmp_2_fu_250_p3 & tmp_1_fu_236_p3);

assign and_ln90_20_fu_2428_p2 = (tmp_45_fu_2254_p3 & tmp_42_fu_2224_p3);

assign and_ln90_21_fu_2718_p2 = (trunc_ln86_9_fu_2516_p1 & tmp_52_fu_2570_p3);

assign and_ln90_22_fu_2724_p2 = (tmp_50_fu_2548_p3 & tmp_49_fu_2534_p3);

assign and_ln90_23_fu_2730_p2 = (tmp_51_fu_2556_p3 & tmp_48_fu_2526_p3);

assign and_ln90_24_fu_3016_p2 = (tmp_60_fu_2868_p3 & tmp_55_fu_2810_p3);

assign and_ln90_25_fu_3022_p2 = (tmp_58_fu_2846_p3 & tmp_57_fu_2832_p3);

assign and_ln90_26_fu_3028_p2 = (tmp_59_fu_2854_p3 & tmp_56_fu_2824_p3);

assign and_ln90_27_fu_3622_p2 = (trunc_ln86_11_fu_3420_p1 & tmp_72_fu_3474_p3);

assign and_ln90_28_fu_3628_p2 = (tmp_70_fu_3452_p3 & tmp_69_fu_3438_p3);

assign and_ln90_29_fu_3634_p2 = (tmp_71_fu_3460_p3 & tmp_68_fu_3430_p3);

assign and_ln90_2_fu_432_p2 = (tmp_fu_228_p3 & tmp_3_fu_258_p3);

assign and_ln90_30_fu_3924_p2 = (trunc_ln86_13_fu_3722_p1 & tmp_78_fu_3776_p3);

assign and_ln90_31_fu_3930_p2 = (tmp_76_fu_3754_p3 & tmp_75_fu_3740_p3);

assign and_ln90_32_fu_3936_p2 = (tmp_77_fu_3762_p3 & tmp_74_fu_3732_p3);

assign and_ln90_33_fu_4222_p2 = (tmp_86_fu_4074_p3 & tmp_81_fu_4016_p3);

assign and_ln90_34_fu_4228_p2 = (tmp_84_fu_4052_p3 & tmp_83_fu_4038_p3);

assign and_ln90_35_fu_4234_p2 = (tmp_85_fu_4060_p3 & tmp_82_fu_4030_p3);

assign and_ln90_36_fu_4626_p2 = (trunc_ln86_15_fu_4424_p1 & tmp_92_fu_4478_p3);

assign and_ln90_37_fu_4632_p2 = (tmp_90_fu_4456_p3 & tmp_89_fu_4442_p3);

assign and_ln90_38_fu_4638_p2 = (tmp_91_fu_4464_p3 & tmp_88_fu_4434_p3);

assign and_ln90_39_fu_4940_p2 = (trunc_ln86_17_fu_4738_p1 & tmp_98_fu_4792_p3);

assign and_ln90_3_fu_722_p2 = (trunc_ln86_3_fu_520_p1 & tmp_10_fu_574_p3);

assign and_ln90_40_fu_4946_p2 = (tmp_96_fu_4770_p3 & tmp_95_fu_4756_p3);

assign and_ln90_41_fu_4952_p2 = (tmp_97_fu_4778_p3 & tmp_94_fu_4748_p3);

assign and_ln90_42_fu_5238_p2 = (tmp_106_fu_5090_p3 & tmp_101_fu_5032_p3);

assign and_ln90_43_fu_5244_p2 = (tmp_104_fu_5068_p3 & tmp_103_fu_5054_p3);

assign and_ln90_44_fu_5250_p2 = (tmp_105_fu_5076_p3 & tmp_102_fu_5046_p3);

assign and_ln90_45_fu_5618_p2 = (tmp_114_fu_5470_p3 & tmp_109_fu_5412_p3);

assign and_ln90_46_fu_5624_p2 = (tmp_112_fu_5448_p3 & tmp_111_fu_5434_p3);

assign and_ln90_47_fu_5630_p2 = (tmp_113_fu_5456_p3 & tmp_110_fu_5426_p3);

assign and_ln90_48_fu_5920_p2 = (trunc_ln86_19_fu_5718_p1 & tmp_120_fu_5772_p3);

assign and_ln90_49_fu_5926_p2 = (tmp_118_fu_5750_p3 & tmp_117_fu_5736_p3);

assign and_ln90_4_fu_728_p2 = (tmp_8_fu_552_p3 & tmp_7_fu_538_p3);

assign and_ln90_50_fu_5932_p2 = (tmp_119_fu_5758_p3 & tmp_116_fu_5728_p3);

assign and_ln90_51_fu_6218_p2 = (tmp_128_fu_6070_p3 & tmp_123_fu_6012_p3);

assign and_ln90_52_fu_6224_p2 = (tmp_126_fu_6048_p3 & tmp_125_fu_6034_p3);

assign and_ln90_53_fu_6230_p2 = (tmp_127_fu_6056_p3 & tmp_124_fu_6026_p3);

assign and_ln90_54_fu_6756_p2 = (tmp_142_fu_6608_p3 & tmp_137_fu_6550_p3);

assign and_ln90_55_fu_6762_p2 = (tmp_140_fu_6586_p3 & tmp_139_fu_6572_p3);

assign and_ln90_56_fu_6768_p2 = (tmp_141_fu_6594_p3 & tmp_138_fu_6564_p3);

assign and_ln90_57_fu_7058_p2 = (trunc_ln86_21_fu_6856_p1 & tmp_148_fu_6910_p3);

assign and_ln90_58_fu_7064_p2 = (tmp_146_fu_6888_p3 & tmp_145_fu_6874_p3);

assign and_ln90_59_fu_7070_p2 = (tmp_147_fu_6896_p3 & tmp_144_fu_6866_p3);

assign and_ln90_5_fu_734_p2 = (tmp_9_fu_560_p3 & tmp_6_fu_530_p3);

assign and_ln90_60_fu_7356_p2 = (tmp_156_fu_7208_p3 & tmp_151_fu_7150_p3);

assign and_ln90_61_fu_7362_p2 = (tmp_154_fu_7186_p3 & tmp_153_fu_7172_p3);

assign and_ln90_62_fu_7368_p2 = (tmp_155_fu_7194_p3 & tmp_152_fu_7164_p3);

assign and_ln90_63_fu_7760_p2 = (trunc_ln86_23_fu_7558_p1 & tmp_162_fu_7612_p3);

assign and_ln90_64_fu_7766_p2 = (tmp_160_fu_7590_p3 & tmp_159_fu_7576_p3);

assign and_ln90_65_fu_7772_p2 = (tmp_161_fu_7598_p3 & tmp_158_fu_7568_p3);

assign and_ln90_66_fu_8074_p2 = (trunc_ln86_25_fu_7872_p1 & tmp_168_fu_7926_p3);

assign and_ln90_67_fu_8080_p2 = (tmp_166_fu_7904_p3 & tmp_165_fu_7890_p3);

assign and_ln90_68_fu_8086_p2 = (tmp_167_fu_7912_p3 & tmp_164_fu_7882_p3);

assign and_ln90_69_fu_8372_p2 = (tmp_176_fu_8224_p3 & tmp_171_fu_8166_p3);

assign and_ln90_6_fu_1020_p2 = (tmp_18_fu_872_p3 & tmp_13_fu_814_p3);

assign and_ln90_70_fu_8378_p2 = (tmp_174_fu_8202_p3 & tmp_173_fu_8188_p3);

assign and_ln90_71_fu_8384_p2 = (tmp_175_fu_8210_p3 & tmp_172_fu_8180_p3);

assign and_ln90_72_fu_8752_p2 = (tmp_184_fu_8604_p3 & tmp_179_fu_8546_p3);

assign and_ln90_73_fu_8758_p2 = (tmp_182_fu_8582_p3 & tmp_181_fu_8568_p3);

assign and_ln90_74_fu_8764_p2 = (tmp_183_fu_8590_p3 & tmp_180_fu_8560_p3);

assign and_ln90_75_fu_9054_p2 = (trunc_ln86_27_fu_8852_p1 & tmp_190_fu_8906_p3);

assign and_ln90_76_fu_9060_p2 = (tmp_188_fu_8884_p3 & tmp_187_fu_8870_p3);

assign and_ln90_77_fu_9066_p2 = (tmp_189_fu_8892_p3 & tmp_186_fu_8862_p3);

assign and_ln90_78_fu_9352_p2 = (tmp_198_fu_9204_p3 & tmp_193_fu_9146_p3);

assign and_ln90_79_fu_9358_p2 = (tmp_196_fu_9182_p3 & tmp_195_fu_9168_p3);

assign and_ln90_7_fu_1026_p2 = (tmp_16_fu_850_p3 & tmp_15_fu_836_p3);

assign and_ln90_80_fu_9364_p2 = (tmp_197_fu_9190_p3 & tmp_194_fu_9160_p3);

assign and_ln90_8_fu_1032_p2 = (tmp_17_fu_858_p3 & tmp_14_fu_828_p3);

assign and_ln90_9_fu_1424_p2 = (trunc_ln86_5_fu_1222_p1 & tmp_24_fu_1276_p3);

assign and_ln90_fu_420_p2 = (trunc_ln86_1_fu_218_p1 & tmp_4_fu_272_p3);

assign and_ln91_10_fu_3942_p2 = (trunc_ln86_12_fu_3718_p1 & tmp_79_fu_3784_p3);

assign and_ln91_11_fu_4240_p2 = (tmp_87_fu_4082_p3 & tmp_80_fu_4008_p3);

assign and_ln91_12_fu_4644_p2 = (trunc_ln86_14_fu_4420_p1 & tmp_93_fu_4486_p3);

assign and_ln91_13_fu_4958_p2 = (trunc_ln86_16_fu_4734_p1 & tmp_99_fu_4800_p3);

assign and_ln91_14_fu_5256_p2 = (tmp_107_fu_5098_p3 & tmp_100_fu_5024_p3);

assign and_ln91_15_fu_5636_p2 = (tmp_115_fu_5478_p3 & tmp_108_fu_5404_p3);

assign and_ln91_16_fu_5938_p2 = (trunc_ln86_18_fu_5714_p1 & tmp_121_fu_5780_p3);

assign and_ln91_17_fu_6236_p2 = (tmp_129_fu_6078_p3 & tmp_122_fu_6004_p3);

assign and_ln91_18_fu_6774_p2 = (tmp_143_fu_6616_p3 & tmp_136_fu_6542_p3);

assign and_ln91_19_fu_7076_p2 = (trunc_ln86_20_fu_6852_p1 & tmp_149_fu_6918_p3);

assign and_ln91_1_fu_740_p2 = (trunc_ln86_2_fu_516_p1 & tmp_11_fu_582_p3);

assign and_ln91_20_fu_7374_p2 = (tmp_157_fu_7216_p3 & tmp_150_fu_7142_p3);

assign and_ln91_21_fu_7778_p2 = (trunc_ln86_22_fu_7554_p1 & tmp_163_fu_7620_p3);

assign and_ln91_22_fu_8092_p2 = (trunc_ln86_24_fu_7868_p1 & tmp_169_fu_7934_p3);

assign and_ln91_23_fu_8390_p2 = (tmp_177_fu_8232_p3 & tmp_170_fu_8158_p3);

assign and_ln91_24_fu_8770_p2 = (tmp_185_fu_8612_p3 & tmp_178_fu_8538_p3);

assign and_ln91_25_fu_9072_p2 = (trunc_ln86_26_fu_8848_p1 & tmp_191_fu_8914_p3);

assign and_ln91_26_fu_9370_p2 = (tmp_199_fu_9212_p3 & tmp_192_fu_9138_p3);

assign and_ln91_2_fu_1038_p2 = (tmp_19_fu_880_p3 & tmp_12_fu_806_p3);

assign and_ln91_3_fu_1442_p2 = (trunc_ln86_4_fu_1218_p1 & tmp_25_fu_1284_p3);

assign and_ln91_4_fu_1756_p2 = (trunc_ln86_6_fu_1532_p1 & tmp_31_fu_1598_p3);

assign and_ln91_5_fu_2054_p2 = (tmp_39_fu_1896_p3 & tmp_32_fu_1822_p3);

assign and_ln91_6_fu_2434_p2 = (tmp_47_fu_2276_p3 & tmp_40_fu_2202_p3);

assign and_ln91_7_fu_2736_p2 = (trunc_ln86_8_fu_2512_p1 & tmp_53_fu_2578_p3);

assign and_ln91_8_fu_3034_p2 = (tmp_61_fu_2876_p3 & tmp_54_fu_2802_p3);

assign and_ln91_9_fu_3640_p2 = (trunc_ln86_10_fu_3416_p1 & tmp_73_fu_3482_p3);

assign and_ln91_fu_438_p2 = (trunc_ln86_fu_214_p1 & tmp_5_fu_280_p3);

assign b0_1_fu_172_p1 = b[7:0];

assign b0_2_fu_200_p1 = b[3:0];

assign b0_3_fu_1182_p4 = {{b[11:8]}};

assign b0_4_fu_3368_p2 = (b0_7_fu_3336_p4 ^ b0_1_fu_172_p1);

assign b0_5_fu_3400_p2 = (b0_8_fu_3326_p4 ^ b0_2_fu_200_p1);

assign b0_6_fu_4384_p4 = {{b_13_fu_3346_p2[11:8]}};

assign b0_7_fu_3336_p4 = {{b[23:16]}};

assign b0_8_fu_3326_p4 = {{b[19:16]}};

assign b0_9_fu_7518_p4 = {{b[27:24]}};

assign b0_fu_144_p1 = b[15:0];

assign b1_11_fu_176_p4 = {{b[15:8]}};

assign b1_12_fu_204_p4 = {{b[7:4]}};

assign b1_13_fu_1208_p4 = {{b_6_fu_1192_p2[7:4]}};

assign b1_14_fu_2192_p4 = {{b[15:12]}};

assign b1_15_fu_3374_p4 = {{b_13_fu_3346_p2[15:8]}};

assign b1_16_fu_3406_p4 = {{b0_4_fu_3368_p2[7:4]}};

assign b1_17_fu_4410_p4 = {{b_18_fu_4394_p2[7:4]}};

assign b1_18_fu_5394_p4 = {{b_13_fu_3346_p2[15:12]}};

assign b1_19_fu_6512_p4 = {{b[31:24]}};

assign b1_20_fu_6532_p4 = {{b[23:20]}};

assign b1_21_fu_7544_p4 = {{b_30_fu_7528_p2[7:4]}};

assign b1_22_fu_8528_p4 = {{b[31:28]}};

assign b1_fu_148_p4 = {{b[31:16]}};

assign b_11_fu_2506_p2 = (b1_14_fu_2192_p4 ^ b0_3_fu_1182_p4);

assign b_13_fu_3346_p2 = (b1_fu_148_p4 ^ b0_fu_144_p1);

assign b_16_fu_3712_p2 = (b1_16_fu_3406_p4 ^ b0_5_fu_3400_p2);

assign b_18_fu_4394_p2 = (b1_15_fu_3374_p4 ^ b0_4_fu_3368_p2);

assign b_19_fu_4728_p2 = (xor_ln99_16_fu_4722_p2 ^ b0_6_fu_4384_p4);

assign b_23_fu_5708_p2 = (b1_18_fu_5394_p4 ^ b0_6_fu_4384_p4);

assign b_28_fu_6846_p2 = (b1_20_fu_6532_p4 ^ b0_8_fu_3326_p4);

assign b_30_fu_7528_p2 = (b1_19_fu_6512_p4 ^ b0_7_fu_3336_p4);

assign b_31_fu_7862_p2 = (xor_ln99_26_fu_7856_p2 ^ b0_8_fu_3326_p4);

assign b_35_fu_8842_p2 = (b1_22_fu_8528_p4 ^ b0_9_fu_7518_p4);

assign b_4_fu_510_p2 = (b1_12_fu_204_p4 ^ b0_2_fu_200_p1);

assign b_6_fu_1192_p2 = (b1_11_fu_176_p4 ^ b0_1_fu_172_p1);

assign b_7_fu_1526_p2 = (xor_ln99_4_fu_1520_p2 ^ b0_3_fu_1182_p4);

assign res_16_fu_4324_p5 = {{{{xor_ln54_7_fu_4318_p2}, {xor_ln53_3_fu_4306_p2}}, {xor_ln91_23_fu_4288_p2}}, {xor_ln88_59_fu_4216_p2}};

assign res_20_fu_5340_p5 = {{{{xor_ln54_9_fu_5334_p2}, {xor_ln53_4_fu_5322_p2}}, {xor_ln91_29_fu_5304_p2}}, {xor_ln88_74_fu_5232_p2}};

assign res_24_fu_6320_p5 = {{{{xor_ln54_11_fu_6314_p2}, {xor_ln53_5_fu_6302_p2}}, {xor_ln91_35_fu_6284_p2}}, {xor_ln88_89_fu_6212_p2}};

assign res_25_fu_6456_p6 = {{{{{xor_ln65_5_fu_6450_p2}, {xor_ln64_3_fu_6416_p2}}, {xor_ln63_1_fu_6392_p2}}, {xor_ln62_1_fu_6370_p2}}, {xor_ln101_25_fu_6344_p2}};

assign res_29_fu_7458_p5 = {{{{xor_ln54_13_fu_7452_p2}, {xor_ln53_6_fu_7440_p2}}, {xor_ln91_41_fu_7422_p2}}, {xor_ln88_104_fu_7350_p2}};

assign res_33_fu_8474_p5 = {{{{xor_ln54_15_fu_8468_p2}, {xor_ln53_7_fu_8456_p2}}, {xor_ln91_47_fu_8438_p2}}, {xor_ln88_119_fu_8366_p2}};

assign res_37_fu_9454_p5 = {{{{xor_ln54_17_fu_9448_p2}, {xor_ln53_8_fu_9436_p2}}, {xor_ln91_53_fu_9418_p2}}, {xor_ln88_134_fu_9346_p2}};

assign res_38_fu_9590_p6 = {{{{{xor_ln65_8_fu_9584_p2}, {xor_ln64_5_fu_9550_p2}}, {xor_ln63_2_fu_9526_p2}}, {xor_ln62_2_fu_9504_p2}}, {xor_ln101_40_fu_9478_p2}};

assign res_39_fu_9742_p6 = {{{{{xor_ln65_11_fu_9726_p2}, {xor_ln64_7_fu_9692_p2}}, {xor_ln63_3_fu_9664_p2}}, {xor_ln62_3_fu_9642_p2}}, {tmp_s_fu_9732_p4}};

assign res_40_fu_492_p5 = {{{{xor_ln91_1_fu_486_p2}, {xor_ln88_4_fu_414_p2}}, {xor_ln87_4_fu_360_p2}}, {xor_ln86_2_fu_306_p2}};

assign res_41_fu_794_p5 = {{{{xor_ln91_3_fu_788_p2}, {xor_ln88_9_fu_716_p2}}, {xor_ln87_9_fu_662_p2}}, {xor_ln86_5_fu_608_p2}};

assign res_42_fu_1092_p5 = {{{{xor_ln91_5_fu_1086_p2}, {xor_ln88_14_fu_1014_p2}}, {xor_ln87_14_fu_960_p2}}, {xor_ln86_8_fu_906_p2}};

assign res_43_fu_1496_p5 = {{{{xor_ln91_7_fu_1490_p2}, {xor_ln88_19_fu_1418_p2}}, {xor_ln87_19_fu_1364_p2}}, {xor_ln86_11_fu_1310_p2}};

assign res_44_fu_1810_p5 = {{{{xor_ln91_9_fu_1804_p2}, {xor_ln88_24_fu_1732_p2}}, {xor_ln87_24_fu_1678_p2}}, {xor_ln86_14_fu_1624_p2}};

assign res_45_fu_2108_p5 = {{{{xor_ln91_11_fu_2102_p2}, {xor_ln88_29_fu_2030_p2}}, {xor_ln87_29_fu_1976_p2}}, {xor_ln86_17_fu_1922_p2}};

assign res_46_fu_2488_p5 = {{{{xor_ln91_13_fu_2482_p2}, {xor_ln88_34_fu_2410_p2}}, {xor_ln87_34_fu_2356_p2}}, {xor_ln86_20_fu_2302_p2}};

assign res_47_fu_2790_p5 = {{{{xor_ln91_15_fu_2784_p2}, {xor_ln88_39_fu_2712_p2}}, {xor_ln87_39_fu_2658_p2}}, {xor_ln86_23_fu_2604_p2}};

assign res_48_fu_3088_p5 = {{{{xor_ln91_17_fu_3082_p2}, {xor_ln88_44_fu_3010_p2}}, {xor_ln87_44_fu_2956_p2}}, {xor_ln86_26_fu_2902_p2}};

assign res_49_fu_3694_p5 = {{{{xor_ln91_19_fu_3688_p2}, {xor_ln88_49_fu_3616_p2}}, {xor_ln87_49_fu_3562_p2}}, {xor_ln86_29_fu_3508_p2}};

assign res_4_fu_2138_p5 = {{{{xor_ln54_3_fu_2132_p2}, {xor_ln53_1_fu_2120_p2}}, {xor_ln91_11_fu_2102_p2}}, {xor_ln88_29_fu_2030_p2}};

assign res_50_fu_3996_p5 = {{{{xor_ln91_21_fu_3990_p2}, {xor_ln88_54_fu_3918_p2}}, {xor_ln87_54_fu_3864_p2}}, {xor_ln86_32_fu_3810_p2}};

assign res_51_fu_4294_p5 = {{{{xor_ln91_23_fu_4288_p2}, {xor_ln88_59_fu_4216_p2}}, {xor_ln87_59_fu_4162_p2}}, {xor_ln86_35_fu_4108_p2}};

assign res_52_fu_4698_p5 = {{{{xor_ln91_25_fu_4692_p2}, {xor_ln88_64_fu_4620_p2}}, {xor_ln87_64_fu_4566_p2}}, {xor_ln86_38_fu_4512_p2}};

assign res_53_fu_5012_p5 = {{{{xor_ln91_27_fu_5006_p2}, {xor_ln88_69_fu_4934_p2}}, {xor_ln87_69_fu_4880_p2}}, {xor_ln86_41_fu_4826_p2}};

assign res_54_fu_5310_p5 = {{{{xor_ln91_29_fu_5304_p2}, {xor_ln88_74_fu_5232_p2}}, {xor_ln87_74_fu_5178_p2}}, {xor_ln86_44_fu_5124_p2}};

assign res_55_fu_5690_p5 = {{{{xor_ln91_31_fu_5684_p2}, {xor_ln88_79_fu_5612_p2}}, {xor_ln87_79_fu_5558_p2}}, {xor_ln86_47_fu_5504_p2}};

assign res_56_fu_5992_p5 = {{{{xor_ln91_33_fu_5986_p2}, {xor_ln88_84_fu_5914_p2}}, {xor_ln87_84_fu_5860_p2}}, {xor_ln86_50_fu_5806_p2}};

assign res_57_fu_6290_p5 = {{{{xor_ln91_35_fu_6284_p2}, {xor_ln88_89_fu_6212_p2}}, {xor_ln87_89_fu_6158_p2}}, {xor_ln86_53_fu_6104_p2}};

assign res_58_fu_6828_p5 = {{{{xor_ln91_37_fu_6822_p2}, {xor_ln88_94_fu_6750_p2}}, {xor_ln87_94_fu_6696_p2}}, {xor_ln86_56_fu_6642_p2}};

assign res_59_fu_7130_p5 = {{{{xor_ln91_39_fu_7124_p2}, {xor_ln88_99_fu_7052_p2}}, {xor_ln87_99_fu_6998_p2}}, {xor_ln86_59_fu_6944_p2}};

assign res_60_fu_7428_p5 = {{{{xor_ln91_41_fu_7422_p2}, {xor_ln88_104_fu_7350_p2}}, {xor_ln87_104_fu_7296_p2}}, {xor_ln86_62_fu_7242_p2}};

assign res_61_fu_7832_p5 = {{{{xor_ln91_43_fu_7826_p2}, {xor_ln88_109_fu_7754_p2}}, {xor_ln87_109_fu_7700_p2}}, {xor_ln86_65_fu_7646_p2}};

assign res_62_fu_8146_p5 = {{{{xor_ln91_45_fu_8140_p2}, {xor_ln88_114_fu_8068_p2}}, {xor_ln87_114_fu_8014_p2}}, {xor_ln86_68_fu_7960_p2}};

assign res_63_fu_8444_p5 = {{{{xor_ln91_47_fu_8438_p2}, {xor_ln88_119_fu_8366_p2}}, {xor_ln87_119_fu_8312_p2}}, {xor_ln86_71_fu_8258_p2}};

assign res_64_fu_8824_p5 = {{{{xor_ln91_49_fu_8818_p2}, {xor_ln88_124_fu_8746_p2}}, {xor_ln87_124_fu_8692_p2}}, {xor_ln86_74_fu_8638_p2}};

assign res_65_fu_9126_p5 = {{{{xor_ln91_51_fu_9120_p2}, {xor_ln88_129_fu_9048_p2}}, {xor_ln87_129_fu_8994_p2}}, {xor_ln86_77_fu_8940_p2}};

assign res_66_fu_9424_p5 = {{{{xor_ln91_53_fu_9418_p2}, {xor_ln88_134_fu_9346_p2}}, {xor_ln87_134_fu_9292_p2}}, {xor_ln86_80_fu_9238_p2}};

assign res_8_fu_3118_p5 = {{{{xor_ln54_5_fu_3112_p2}, {xor_ln53_2_fu_3100_p2}}, {xor_ln91_17_fu_3082_p2}}, {xor_ln88_44_fu_3010_p2}};

assign res_9_fu_3254_p6 = {{{{{xor_ln65_2_fu_3248_p2}, {xor_ln64_1_fu_3214_p2}}, {xor_ln63_fu_3190_p2}}, {xor_ln62_fu_3168_p2}}, {xor_ln101_10_fu_3142_p2}};

assign res_fu_1122_p5 = {{{{xor_ln54_1_fu_1116_p2}, {xor_ln53_fu_1104_p2}}, {xor_ln91_5_fu_1086_p2}}, {xor_ln88_14_fu_1014_p2}};

assign tmp_100_fu_5024_p3 = a_23_fu_4378_p2[32'd4];

assign tmp_101_fu_5032_p3 = b_18_fu_4394_p2[32'd4];

assign tmp_102_fu_5046_p3 = a_23_fu_4378_p2[32'd5];

assign tmp_103_fu_5054_p3 = b_18_fu_4394_p2[32'd5];

assign tmp_104_fu_5068_p3 = a_23_fu_4378_p2[32'd6];

assign tmp_105_fu_5076_p3 = b_18_fu_4394_p2[32'd6];

assign tmp_106_fu_5090_p3 = a_23_fu_4378_p2[32'd7];

assign tmp_107_fu_5098_p3 = b_18_fu_4394_p2[32'd7];

assign tmp_108_fu_5404_p3 = a_17_fu_3320_p2[32'd8];

assign tmp_109_fu_5412_p3 = b_13_fu_3346_p2[32'd8];

assign tmp_10_fu_574_p3 = a_4_fu_504_p2[32'd3];

assign tmp_110_fu_5426_p3 = a_17_fu_3320_p2[32'd9];

assign tmp_111_fu_5434_p3 = b_13_fu_3346_p2[32'd9];

assign tmp_112_fu_5448_p3 = a_17_fu_3320_p2[32'd10];

assign tmp_113_fu_5456_p3 = b_13_fu_3346_p2[32'd10];

assign tmp_114_fu_5470_p3 = a_17_fu_3320_p2[32'd11];

assign tmp_115_fu_5478_p3 = b_13_fu_3346_p2[32'd11];

assign tmp_116_fu_5728_p3 = a_29_fu_5702_p2[32'd1];

assign tmp_117_fu_5736_p3 = b_23_fu_5708_p2[32'd1];

assign tmp_118_fu_5750_p3 = a_29_fu_5702_p2[32'd2];

assign tmp_119_fu_5758_p3 = b_23_fu_5708_p2[32'd2];

assign tmp_11_fu_582_p3 = b_4_fu_510_p2[32'd3];

assign tmp_120_fu_5772_p3 = a_29_fu_5702_p2[32'd3];

assign tmp_121_fu_5780_p3 = b_23_fu_5708_p2[32'd3];

assign tmp_122_fu_6004_p3 = a_17_fu_3320_p2[32'd12];

assign tmp_123_fu_6012_p3 = b_13_fu_3346_p2[32'd12];

assign tmp_124_fu_6026_p3 = a_17_fu_3320_p2[32'd13];

assign tmp_125_fu_6034_p3 = b_13_fu_3346_p2[32'd13];

assign tmp_126_fu_6048_p3 = a_17_fu_3320_p2[32'd14];

assign tmp_127_fu_6056_p3 = b_13_fu_3346_p2[32'd14];

assign tmp_128_fu_6070_p3 = a_17_fu_3320_p2[32'd15];

assign tmp_129_fu_6078_p3 = b_13_fu_3346_p2[32'd15];

assign tmp_12_fu_806_p3 = a[32'd4];

assign tmp_130_fu_6362_p3 = xor_ln101_25_fu_6344_p2[32'd2];

assign tmp_131_fu_6376_p3 = xor_ln101_23_fu_6332_p2[32'd1];

assign tmp_132_fu_6384_p3 = xor_ln101_25_fu_6344_p2[32'd3];

assign tmp_133_fu_6398_p3 = xor_ln101_23_fu_6332_p2[32'd2];

assign tmp_134_fu_6422_p3 = xor_ln101_23_fu_6332_p2[32'd3];

assign tmp_135_fu_6430_p3 = xor_ln101_25_fu_6344_p2[32'd1];

assign tmp_136_fu_6542_p3 = a[32'd16];

assign tmp_137_fu_6550_p3 = b[32'd16];

assign tmp_138_fu_6564_p3 = a[32'd17];

assign tmp_139_fu_6572_p3 = b[32'd17];

assign tmp_13_fu_814_p3 = b[32'd4];

assign tmp_140_fu_6586_p3 = a[32'd18];

assign tmp_141_fu_6594_p3 = b[32'd18];

assign tmp_142_fu_6608_p3 = a[32'd19];

assign tmp_143_fu_6616_p3 = b[32'd19];

assign tmp_144_fu_6866_p3 = a_36_fu_6840_p2[32'd1];

assign tmp_145_fu_6874_p3 = b_28_fu_6846_p2[32'd1];

assign tmp_146_fu_6888_p3 = a_36_fu_6840_p2[32'd2];

assign tmp_147_fu_6896_p3 = b_28_fu_6846_p2[32'd2];

assign tmp_148_fu_6910_p3 = a_36_fu_6840_p2[32'd3];

assign tmp_149_fu_6918_p3 = b_28_fu_6846_p2[32'd3];

assign tmp_14_fu_828_p3 = a[32'd5];

assign tmp_150_fu_7142_p3 = a[32'd20];

assign tmp_151_fu_7150_p3 = b[32'd20];

assign tmp_152_fu_7164_p3 = a[32'd21];

assign tmp_153_fu_7172_p3 = b[32'd21];

assign tmp_154_fu_7186_p3 = a[32'd22];

assign tmp_155_fu_7194_p3 = b[32'd22];

assign tmp_156_fu_7208_p3 = a[32'd23];

assign tmp_157_fu_7216_p3 = b[32'd23];

assign tmp_158_fu_7568_p3 = a_39_fu_7512_p2[32'd1];

assign tmp_159_fu_7576_p3 = b_30_fu_7528_p2[32'd1];

assign tmp_15_fu_836_p3 = b[32'd5];

assign tmp_160_fu_7590_p3 = a_39_fu_7512_p2[32'd2];

assign tmp_161_fu_7598_p3 = b_30_fu_7528_p2[32'd2];

assign tmp_162_fu_7612_p3 = a_39_fu_7512_p2[32'd3];

assign tmp_163_fu_7620_p3 = b_30_fu_7528_p2[32'd3];

assign tmp_164_fu_7882_p3 = a_40_fu_7850_p2[32'd1];

assign tmp_165_fu_7890_p3 = b_31_fu_7862_p2[32'd1];

assign tmp_166_fu_7904_p3 = a_40_fu_7850_p2[32'd2];

assign tmp_167_fu_7912_p3 = b_31_fu_7862_p2[32'd2];

assign tmp_168_fu_7926_p3 = a_40_fu_7850_p2[32'd3];

assign tmp_169_fu_7934_p3 = b_31_fu_7862_p2[32'd3];

assign tmp_16_fu_850_p3 = a[32'd6];

assign tmp_170_fu_8158_p3 = a_39_fu_7512_p2[32'd4];

assign tmp_171_fu_8166_p3 = b_30_fu_7528_p2[32'd4];

assign tmp_172_fu_8180_p3 = a_39_fu_7512_p2[32'd5];

assign tmp_173_fu_8188_p3 = b_30_fu_7528_p2[32'd5];

assign tmp_174_fu_8202_p3 = a_39_fu_7512_p2[32'd6];

assign tmp_175_fu_8210_p3 = b_30_fu_7528_p2[32'd6];

assign tmp_176_fu_8224_p3 = a_39_fu_7512_p2[32'd7];

assign tmp_177_fu_8232_p3 = b_30_fu_7528_p2[32'd7];

assign tmp_178_fu_8538_p3 = a[32'd24];

assign tmp_179_fu_8546_p3 = b[32'd24];

assign tmp_17_fu_858_p3 = b[32'd6];

assign tmp_180_fu_8560_p3 = a[32'd25];

assign tmp_181_fu_8568_p3 = b[32'd25];

assign tmp_182_fu_8582_p3 = a[32'd26];

assign tmp_183_fu_8590_p3 = b[32'd26];

assign tmp_184_fu_8604_p3 = a[32'd27];

assign tmp_185_fu_8612_p3 = b[32'd27];

assign tmp_186_fu_8862_p3 = a_45_fu_8836_p2[32'd1];

assign tmp_187_fu_8870_p3 = b_35_fu_8842_p2[32'd1];

assign tmp_188_fu_8884_p3 = a_45_fu_8836_p2[32'd2];

assign tmp_189_fu_8892_p3 = b_35_fu_8842_p2[32'd2];

assign tmp_18_fu_872_p3 = a[32'd7];

assign tmp_190_fu_8906_p3 = a_45_fu_8836_p2[32'd3];

assign tmp_191_fu_8914_p3 = b_35_fu_8842_p2[32'd3];

assign tmp_192_fu_9138_p3 = a[32'd28];

assign tmp_193_fu_9146_p3 = b[32'd28];

assign tmp_194_fu_9160_p3 = a[32'd29];

assign tmp_195_fu_9168_p3 = b[32'd29];

assign tmp_196_fu_9182_p3 = a[32'd30];

assign tmp_197_fu_9190_p3 = b[32'd30];

assign tmp_198_fu_9204_p3 = a[32'd31];

assign tmp_199_fu_9212_p3 = b[32'd31];

assign tmp_19_fu_880_p3 = b[32'd7];

assign tmp_1_fu_236_p3 = b[32'd1];

assign tmp_200_fu_9496_p3 = xor_ln101_40_fu_9478_p2[32'd2];

assign tmp_201_fu_9510_p3 = xor_ln101_38_fu_9466_p2[32'd1];

assign tmp_202_fu_9518_p3 = xor_ln101_40_fu_9478_p2[32'd3];

assign tmp_203_fu_9532_p3 = xor_ln101_38_fu_9466_p2[32'd2];

assign tmp_204_fu_9556_p3 = xor_ln101_38_fu_9466_p2[32'd3];

assign tmp_205_fu_9564_p3 = xor_ln101_40_fu_9478_p2[32'd1];

assign tmp_206_fu_9634_p3 = a1_23_fu_9616_p2[32'd6];

assign tmp_207_fu_9648_p3 = a1_23_fu_9616_p2[32'd1];

assign tmp_208_fu_9656_p3 = a1_23_fu_9616_p2[32'd7];

assign tmp_209_fu_9670_p3 = a1_23_fu_9616_p2[32'd2];

assign tmp_20_fu_1232_p3 = a_7_fu_1176_p2[32'd1];

assign tmp_210_fu_9678_p3 = a1_23_fu_9616_p2[32'd4];

assign tmp_211_fu_9698_p3 = a1_23_fu_9616_p2[32'd3];

assign tmp_212_fu_9706_p3 = a1_23_fu_9616_p2[32'd5];

assign tmp_213_fu_9762_p3 = {{xor_ln70_fu_9756_p2}, {a1_23_fu_9616_p2}};

assign tmp_21_fu_1240_p3 = b_6_fu_1192_p2[32'd1];

assign tmp_22_fu_1254_p3 = a_7_fu_1176_p2[32'd2];

assign tmp_23_fu_1262_p3 = b_6_fu_1192_p2[32'd2];

assign tmp_24_fu_1276_p3 = a_7_fu_1176_p2[32'd3];

assign tmp_25_fu_1284_p3 = b_6_fu_1192_p2[32'd3];

assign tmp_26_fu_1546_p3 = a_8_fu_1514_p2[32'd1];

assign tmp_27_fu_1554_p3 = b_7_fu_1526_p2[32'd1];

assign tmp_28_fu_1568_p3 = a_8_fu_1514_p2[32'd2];

assign tmp_29_fu_1576_p3 = b_7_fu_1526_p2[32'd2];

assign tmp_2_fu_250_p3 = a[32'd2];

assign tmp_30_fu_1590_p3 = a_8_fu_1514_p2[32'd3];

assign tmp_31_fu_1598_p3 = b_7_fu_1526_p2[32'd3];

assign tmp_32_fu_1822_p3 = a_7_fu_1176_p2[32'd4];

assign tmp_33_fu_1830_p3 = b_6_fu_1192_p2[32'd4];

assign tmp_34_fu_1844_p3 = a_7_fu_1176_p2[32'd5];

assign tmp_35_fu_1852_p3 = b_6_fu_1192_p2[32'd5];

assign tmp_36_fu_1866_p3 = a_7_fu_1176_p2[32'd6];

assign tmp_37_fu_1874_p3 = b_6_fu_1192_p2[32'd6];

assign tmp_38_fu_1888_p3 = a_7_fu_1176_p2[32'd7];

assign tmp_39_fu_1896_p3 = b_6_fu_1192_p2[32'd7];

assign tmp_3_fu_258_p3 = b[32'd2];

assign tmp_40_fu_2202_p3 = a[32'd8];

assign tmp_41_fu_2210_p3 = b[32'd8];

assign tmp_42_fu_2224_p3 = a[32'd9];

assign tmp_43_fu_2232_p3 = b[32'd9];

assign tmp_44_fu_2246_p3 = a[32'd10];

assign tmp_45_fu_2254_p3 = b[32'd10];

assign tmp_46_fu_2268_p3 = a[32'd11];

assign tmp_47_fu_2276_p3 = b[32'd11];

assign tmp_48_fu_2526_p3 = a_13_fu_2500_p2[32'd1];

assign tmp_49_fu_2534_p3 = b_11_fu_2506_p2[32'd1];

assign tmp_4_fu_272_p3 = a[32'd3];

assign tmp_50_fu_2548_p3 = a_13_fu_2500_p2[32'd2];

assign tmp_51_fu_2556_p3 = b_11_fu_2506_p2[32'd2];

assign tmp_52_fu_2570_p3 = a_13_fu_2500_p2[32'd3];

assign tmp_53_fu_2578_p3 = b_11_fu_2506_p2[32'd3];

assign tmp_54_fu_2802_p3 = a[32'd12];

assign tmp_55_fu_2810_p3 = b[32'd12];

assign tmp_56_fu_2824_p3 = a[32'd13];

assign tmp_57_fu_2832_p3 = b[32'd13];

assign tmp_58_fu_2846_p3 = a[32'd14];

assign tmp_59_fu_2854_p3 = b[32'd14];

assign tmp_5_fu_280_p3 = b[32'd3];

assign tmp_60_fu_2868_p3 = a[32'd15];

assign tmp_61_fu_2876_p3 = b[32'd15];

assign tmp_62_fu_3160_p3 = xor_ln101_10_fu_3142_p2[32'd2];

assign tmp_63_fu_3174_p3 = xor_ln101_8_fu_3130_p2[32'd1];

assign tmp_64_fu_3182_p3 = xor_ln101_10_fu_3142_p2[32'd3];

assign tmp_65_fu_3196_p3 = xor_ln101_8_fu_3130_p2[32'd2];

assign tmp_66_fu_3220_p3 = xor_ln101_8_fu_3130_p2[32'd3];

assign tmp_67_fu_3228_p3 = xor_ln101_10_fu_3142_p2[32'd1];

assign tmp_68_fu_3430_p3 = a_17_fu_3320_p2[32'd1];

assign tmp_69_fu_3438_p3 = b_13_fu_3346_p2[32'd1];

assign tmp_6_fu_530_p3 = a_4_fu_504_p2[32'd1];

assign tmp_70_fu_3452_p3 = a_17_fu_3320_p2[32'd2];

assign tmp_71_fu_3460_p3 = b_13_fu_3346_p2[32'd2];

assign tmp_72_fu_3474_p3 = a_17_fu_3320_p2[32'd3];

assign tmp_73_fu_3482_p3 = b_13_fu_3346_p2[32'd3];

assign tmp_74_fu_3732_p3 = a_20_fu_3706_p2[32'd1];

assign tmp_75_fu_3740_p3 = b_16_fu_3712_p2[32'd1];

assign tmp_76_fu_3754_p3 = a_20_fu_3706_p2[32'd2];

assign tmp_77_fu_3762_p3 = b_16_fu_3712_p2[32'd2];

assign tmp_78_fu_3776_p3 = a_20_fu_3706_p2[32'd3];

assign tmp_79_fu_3784_p3 = b_16_fu_3712_p2[32'd3];

assign tmp_7_fu_538_p3 = b_4_fu_510_p2[32'd1];

assign tmp_80_fu_4008_p3 = a0_15_fu_3352_p2[32'd4];

assign tmp_81_fu_4016_p3 = b0_4_fu_3368_p2[32'd4];

assign tmp_82_fu_4030_p3 = a0_15_fu_3352_p2[32'd5];

assign tmp_83_fu_4038_p3 = b0_4_fu_3368_p2[32'd5];

assign tmp_84_fu_4052_p3 = a0_15_fu_3352_p2[32'd6];

assign tmp_85_fu_4060_p3 = b0_4_fu_3368_p2[32'd6];

assign tmp_86_fu_4074_p3 = a0_15_fu_3352_p2[32'd7];

assign tmp_87_fu_4082_p3 = b0_4_fu_3368_p2[32'd7];

assign tmp_88_fu_4434_p3 = a_23_fu_4378_p2[32'd1];

assign tmp_89_fu_4442_p3 = b_18_fu_4394_p2[32'd1];

assign tmp_8_fu_552_p3 = a_4_fu_504_p2[32'd2];

assign tmp_90_fu_4456_p3 = a_23_fu_4378_p2[32'd2];

assign tmp_91_fu_4464_p3 = b_18_fu_4394_p2[32'd2];

assign tmp_92_fu_4478_p3 = a_23_fu_4378_p2[32'd3];

assign tmp_93_fu_4486_p3 = b_18_fu_4394_p2[32'd3];

assign tmp_94_fu_4748_p3 = a_24_fu_4716_p2[32'd1];

assign tmp_95_fu_4756_p3 = b_19_fu_4728_p2[32'd1];

assign tmp_96_fu_4770_p3 = a_24_fu_4716_p2[32'd2];

assign tmp_97_fu_4778_p3 = b_19_fu_4728_p2[32'd2];

assign tmp_98_fu_4792_p3 = a_24_fu_4716_p2[32'd3];

assign tmp_99_fu_4800_p3 = b_19_fu_4728_p2[32'd3];

assign tmp_9_fu_560_p3 = b_4_fu_510_p2[32'd2];

assign tmp_fu_228_p3 = a[32'd1];

assign tmp_s_fu_9732_p4 = {{a1_23_fu_9616_p2[7:4]}};

assign trunc_ln62_1_fu_6358_p1 = xor_ln101_23_fu_6332_p2[0:0];

assign trunc_ln62_2_fu_9492_p1 = xor_ln101_38_fu_9466_p2[0:0];

assign trunc_ln62_3_fu_9630_p1 = a1_23_fu_9616_p2[0:0];

assign trunc_ln62_fu_3156_p1 = xor_ln101_8_fu_3130_p2[0:0];

assign trunc_ln64_1_fu_6406_p1 = xor_ln101_25_fu_6344_p2[0:0];

assign trunc_ln64_2_fu_9540_p1 = xor_ln101_40_fu_9478_p2[0:0];

assign trunc_ln64_fu_3204_p1 = xor_ln101_10_fu_3142_p2[0:0];

assign trunc_ln86_10_fu_3416_p1 = a_17_fu_3320_p2[0:0];

assign trunc_ln86_11_fu_3420_p1 = b_13_fu_3346_p2[0:0];

assign trunc_ln86_12_fu_3718_p1 = a_20_fu_3706_p2[0:0];

assign trunc_ln86_13_fu_3722_p1 = b_16_fu_3712_p2[0:0];

assign trunc_ln86_14_fu_4420_p1 = a_23_fu_4378_p2[0:0];

assign trunc_ln86_15_fu_4424_p1 = b_18_fu_4394_p2[0:0];

assign trunc_ln86_16_fu_4734_p1 = a_24_fu_4716_p2[0:0];

assign trunc_ln86_17_fu_4738_p1 = b_19_fu_4728_p2[0:0];

assign trunc_ln86_18_fu_5714_p1 = a_29_fu_5702_p2[0:0];

assign trunc_ln86_19_fu_5718_p1 = b_23_fu_5708_p2[0:0];

assign trunc_ln86_1_fu_218_p1 = b[0:0];

assign trunc_ln86_20_fu_6852_p1 = a_36_fu_6840_p2[0:0];

assign trunc_ln86_21_fu_6856_p1 = b_28_fu_6846_p2[0:0];

assign trunc_ln86_22_fu_7554_p1 = a_39_fu_7512_p2[0:0];

assign trunc_ln86_23_fu_7558_p1 = b_30_fu_7528_p2[0:0];

assign trunc_ln86_24_fu_7868_p1 = a_40_fu_7850_p2[0:0];

assign trunc_ln86_25_fu_7872_p1 = b_31_fu_7862_p2[0:0];

assign trunc_ln86_26_fu_8848_p1 = a_45_fu_8836_p2[0:0];

assign trunc_ln86_27_fu_8852_p1 = b_35_fu_8842_p2[0:0];

assign trunc_ln86_2_fu_516_p1 = a_4_fu_504_p2[0:0];

assign trunc_ln86_3_fu_520_p1 = b_4_fu_510_p2[0:0];

assign trunc_ln86_4_fu_1218_p1 = a_7_fu_1176_p2[0:0];

assign trunc_ln86_5_fu_1222_p1 = b_6_fu_1192_p2[0:0];

assign trunc_ln86_6_fu_1532_p1 = a_8_fu_1514_p2[0:0];

assign trunc_ln86_7_fu_1536_p1 = b_7_fu_1526_p2[0:0];

assign trunc_ln86_8_fu_2512_p1 = a_13_fu_2500_p2[0:0];

assign trunc_ln86_9_fu_2516_p1 = b_11_fu_2506_p2[0:0];

assign trunc_ln86_fu_214_p1 = a[0:0];

assign xor_ln101_10_fu_3142_p2 = (xor_ln101_9_fu_3136_p2 ^ xor_ln101_8_fu_3130_p2);

assign xor_ln101_11_fu_3268_p2 = (z1_2_fu_2174_p3 ^ z0_1_fu_1158_p3);

assign xor_ln101_12_fu_3274_p2 = (z2_fu_3148_p3 ^ res_9_fu_3254_p6);

assign xor_ln101_13_fu_3280_p2 = (xor_ln101_12_fu_3274_p2 ^ xor_ln101_11_fu_3268_p2);

assign xor_ln101_14_fu_3286_p2 = (z2_fu_3148_p3 ^ z0_1_fu_1158_p3);

assign xor_ln101_15_fu_4336_p2 = (res_50_fu_3996_p5 ^ res_49_fu_3694_p5);

assign xor_ln101_16_fu_4342_p2 = (res_51_fu_4294_p5 ^ res_16_fu_4324_p5);

assign xor_ln101_17_fu_4348_p2 = (xor_ln101_16_fu_4342_p2 ^ xor_ln101_15_fu_4336_p2);

assign xor_ln101_18_fu_4354_p2 = (res_51_fu_4294_p5 ^ res_49_fu_3694_p5);

assign xor_ln101_19_fu_5352_p2 = (res_53_fu_5012_p5 ^ res_52_fu_4698_p5);

assign xor_ln101_1_fu_1140_p2 = (res_fu_1122_p5 ^ res_42_fu_1092_p5);

assign xor_ln101_20_fu_5358_p2 = (res_54_fu_5310_p5 ^ res_20_fu_5340_p5);

assign xor_ln101_21_fu_5364_p2 = (xor_ln101_20_fu_5358_p2 ^ xor_ln101_19_fu_5352_p2);

assign xor_ln101_22_fu_5370_p2 = (res_54_fu_5310_p5 ^ res_52_fu_4698_p5);

assign xor_ln101_23_fu_6332_p2 = (res_57_fu_6290_p5 ^ res_55_fu_5690_p5);

assign xor_ln101_24_fu_6338_p2 = (res_56_fu_5992_p5 ^ res_24_fu_6320_p5);

assign xor_ln101_25_fu_6344_p2 = (xor_ln101_24_fu_6338_p2 ^ xor_ln101_23_fu_6332_p2);

assign xor_ln101_26_fu_6470_p2 = (z1_6_fu_5376_p3 ^ z0_6_fu_4360_p3);

assign xor_ln101_27_fu_6476_p2 = (z2_4_fu_6350_p3 ^ res_25_fu_6456_p6);

assign xor_ln101_28_fu_6482_p2 = (xor_ln101_27_fu_6476_p2 ^ xor_ln101_26_fu_6470_p2);

assign xor_ln101_29_fu_6488_p2 = (z2_4_fu_6350_p3 ^ z0_6_fu_4360_p3);

assign xor_ln101_2_fu_1146_p2 = (xor_ln101_fu_1134_p2 ^ xor_ln101_1_fu_1140_p2);

assign xor_ln101_30_fu_7470_p2 = (res_59_fu_7130_p5 ^ res_58_fu_6828_p5);

assign xor_ln101_31_fu_7476_p2 = (res_60_fu_7428_p5 ^ res_29_fu_7458_p5);

assign xor_ln101_32_fu_7482_p2 = (xor_ln101_31_fu_7476_p2 ^ xor_ln101_30_fu_7470_p2);

assign xor_ln101_33_fu_7488_p2 = (res_60_fu_7428_p5 ^ res_58_fu_6828_p5);

assign xor_ln101_34_fu_8486_p2 = (res_62_fu_8146_p5 ^ res_61_fu_7832_p5);

assign xor_ln101_35_fu_8492_p2 = (res_63_fu_8444_p5 ^ res_33_fu_8474_p5);

assign xor_ln101_36_fu_8498_p2 = (xor_ln101_35_fu_8492_p2 ^ xor_ln101_34_fu_8486_p2);

assign xor_ln101_37_fu_8504_p2 = (res_63_fu_8444_p5 ^ res_61_fu_7832_p5);

assign xor_ln101_38_fu_9466_p2 = (res_66_fu_9424_p5 ^ res_64_fu_8824_p5);

assign xor_ln101_39_fu_9472_p2 = (res_65_fu_9126_p5 ^ res_37_fu_9454_p5);

assign xor_ln101_3_fu_1152_p2 = (res_42_fu_1092_p5 ^ res_40_fu_492_p5);

assign xor_ln101_40_fu_9478_p2 = (xor_ln101_39_fu_9472_p2 ^ xor_ln101_38_fu_9466_p2);

assign xor_ln101_42_fu_9610_p2 = (z1_11_fu_8510_p3 ^ res_38_fu_9590_p6);

assign xor_ln101_44_fu_9770_p2 = (z1_8_fu_6494_p3 ^ z0_4_fu_3292_p3);

assign xor_ln101_45_fu_9776_p2 = (z2_6_fu_9622_p3 ^ tmp_213_fu_9762_p3);

assign xor_ln101_46_fu_9782_p2 = (xor_ln101_45_fu_9776_p2 ^ xor_ln101_44_fu_9770_p2);

assign xor_ln101_47_fu_9788_p2 = (z2_6_fu_9622_p3 ^ z0_4_fu_3292_p3);

assign xor_ln101_4_fu_2150_p2 = (res_44_fu_1810_p5 ^ res_43_fu_1496_p5);

assign xor_ln101_5_fu_2156_p2 = (res_4_fu_2138_p5 ^ res_45_fu_2108_p5);

assign xor_ln101_6_fu_2162_p2 = (xor_ln101_5_fu_2156_p2 ^ xor_ln101_4_fu_2150_p2);

assign xor_ln101_7_fu_2168_p2 = (res_45_fu_2108_p5 ^ res_43_fu_1496_p5);

assign xor_ln101_8_fu_3130_p2 = (res_48_fu_3088_p5 ^ res_46_fu_2488_p5);

assign xor_ln101_9_fu_3136_p2 = (res_8_fu_3118_p5 ^ res_47_fu_2790_p5);

assign xor_ln101_fu_1134_p2 = (res_41_fu_794_p5 ^ res_40_fu_492_p5);

assign xor_ln53_1_fu_2120_p2 = (xor_ln91_11_fu_2102_p2 ^ xor_ln86_17_fu_1922_p2);

assign xor_ln53_2_fu_3100_p2 = (xor_ln91_17_fu_3082_p2 ^ xor_ln86_26_fu_2902_p2);

assign xor_ln53_3_fu_4306_p2 = (xor_ln91_23_fu_4288_p2 ^ xor_ln86_35_fu_4108_p2);

assign xor_ln53_4_fu_5322_p2 = (xor_ln91_29_fu_5304_p2 ^ xor_ln86_44_fu_5124_p2);

assign xor_ln53_5_fu_6302_p2 = (xor_ln91_35_fu_6284_p2 ^ xor_ln86_53_fu_6104_p2);

assign xor_ln53_6_fu_7440_p2 = (xor_ln91_41_fu_7422_p2 ^ xor_ln86_62_fu_7242_p2);

assign xor_ln53_7_fu_8456_p2 = (xor_ln91_47_fu_8438_p2 ^ xor_ln86_71_fu_8258_p2);

assign xor_ln53_8_fu_9436_p2 = (xor_ln91_53_fu_9418_p2 ^ xor_ln86_80_fu_9238_p2);

assign xor_ln53_fu_1104_p2 = (xor_ln91_5_fu_1086_p2 ^ xor_ln86_8_fu_906_p2);

assign xor_ln54_10_fu_6308_p2 = (xor_ln91_35_fu_6284_p2 ^ xor_ln88_88_fu_6206_p2);

assign xor_ln54_11_fu_6314_p2 = (xor_ln87_87_fu_6140_p2 ^ xor_ln54_10_fu_6308_p2);

assign xor_ln54_12_fu_7446_p2 = (xor_ln91_41_fu_7422_p2 ^ xor_ln88_103_fu_7344_p2);

assign xor_ln54_13_fu_7452_p2 = (xor_ln87_102_fu_7278_p2 ^ xor_ln54_12_fu_7446_p2);

assign xor_ln54_14_fu_8462_p2 = (xor_ln91_47_fu_8438_p2 ^ xor_ln88_118_fu_8360_p2);

assign xor_ln54_15_fu_8468_p2 = (xor_ln87_117_fu_8294_p2 ^ xor_ln54_14_fu_8462_p2);

assign xor_ln54_16_fu_9442_p2 = (xor_ln91_53_fu_9418_p2 ^ xor_ln88_133_fu_9340_p2);

assign xor_ln54_17_fu_9448_p2 = (xor_ln87_132_fu_9274_p2 ^ xor_ln54_16_fu_9442_p2);

assign xor_ln54_1_fu_1116_p2 = (xor_ln87_12_fu_942_p2 ^ xor_ln54_fu_1110_p2);

assign xor_ln54_2_fu_2126_p2 = (xor_ln91_11_fu_2102_p2 ^ xor_ln88_28_fu_2024_p2);

assign xor_ln54_3_fu_2132_p2 = (xor_ln87_27_fu_1958_p2 ^ xor_ln54_2_fu_2126_p2);

assign xor_ln54_4_fu_3106_p2 = (xor_ln91_17_fu_3082_p2 ^ xor_ln88_43_fu_3004_p2);

assign xor_ln54_5_fu_3112_p2 = (xor_ln87_42_fu_2938_p2 ^ xor_ln54_4_fu_3106_p2);

assign xor_ln54_6_fu_4312_p2 = (xor_ln91_23_fu_4288_p2 ^ xor_ln88_58_fu_4210_p2);

assign xor_ln54_7_fu_4318_p2 = (xor_ln87_57_fu_4144_p2 ^ xor_ln54_6_fu_4312_p2);

assign xor_ln54_8_fu_5328_p2 = (xor_ln91_29_fu_5304_p2 ^ xor_ln88_73_fu_5226_p2);

assign xor_ln54_9_fu_5334_p2 = (xor_ln87_72_fu_5160_p2 ^ xor_ln54_8_fu_5328_p2);

assign xor_ln54_fu_1110_p2 = (xor_ln91_5_fu_1086_p2 ^ xor_ln88_13_fu_1008_p2);

assign xor_ln62_1_fu_6370_p2 = (trunc_ln62_1_fu_6358_p1 ^ tmp_130_fu_6362_p3);

assign xor_ln62_2_fu_9504_p2 = (trunc_ln62_2_fu_9492_p1 ^ tmp_200_fu_9496_p3);

assign xor_ln62_3_fu_9642_p2 = (trunc_ln62_3_fu_9630_p1 ^ tmp_206_fu_9634_p3);

assign xor_ln62_fu_3168_p2 = (trunc_ln62_fu_3156_p1 ^ tmp_62_fu_3160_p3);

assign xor_ln63_1_fu_6392_p2 = (tmp_132_fu_6384_p3 ^ tmp_131_fu_6376_p3);

assign xor_ln63_2_fu_9526_p2 = (tmp_202_fu_9518_p3 ^ tmp_201_fu_9510_p3);

assign xor_ln63_3_fu_9664_p2 = (tmp_208_fu_9656_p3 ^ tmp_207_fu_9648_p3);

assign xor_ln63_fu_3190_p2 = (tmp_64_fu_3182_p3 ^ tmp_63_fu_3174_p3);

assign xor_ln64_1_fu_3214_p2 = (xor_ln64_fu_3208_p2 ^ tmp_65_fu_3196_p3);

assign xor_ln64_2_fu_6410_p2 = (trunc_ln64_1_fu_6406_p1 ^ tmp_132_fu_6384_p3);

assign xor_ln64_3_fu_6416_p2 = (xor_ln64_2_fu_6410_p2 ^ tmp_133_fu_6398_p3);

assign xor_ln64_4_fu_9544_p2 = (trunc_ln64_2_fu_9540_p1 ^ tmp_202_fu_9518_p3);

assign xor_ln64_5_fu_9550_p2 = (xor_ln64_4_fu_9544_p2 ^ tmp_203_fu_9532_p3);

assign xor_ln64_6_fu_9686_p2 = (tmp_210_fu_9678_p3 ^ tmp_208_fu_9656_p3);

assign xor_ln64_7_fu_9692_p2 = (xor_ln64_6_fu_9686_p2 ^ tmp_209_fu_9670_p3);

assign xor_ln64_fu_3208_p2 = (trunc_ln64_fu_3204_p1 ^ tmp_64_fu_3182_p3);

assign xor_ln65_10_fu_9720_p2 = (tmp_208_fu_9656_p3 ^ tmp_206_fu_9634_p3);

assign xor_ln65_11_fu_9726_p2 = (xor_ln65_9_fu_9714_p2 ^ xor_ln65_10_fu_9720_p2);

assign xor_ln65_1_fu_3242_p2 = (tmp_64_fu_3182_p3 ^ tmp_62_fu_3160_p3);

assign xor_ln65_2_fu_3248_p2 = (xor_ln65_fu_3236_p2 ^ xor_ln65_1_fu_3242_p2);

assign xor_ln65_3_fu_6438_p2 = (tmp_135_fu_6430_p3 ^ tmp_134_fu_6422_p3);

assign xor_ln65_4_fu_6444_p2 = (tmp_132_fu_6384_p3 ^ tmp_130_fu_6362_p3);

assign xor_ln65_5_fu_6450_p2 = (xor_ln65_4_fu_6444_p2 ^ xor_ln65_3_fu_6438_p2);

assign xor_ln65_6_fu_9572_p2 = (tmp_205_fu_9564_p3 ^ tmp_204_fu_9556_p3);

assign xor_ln65_7_fu_9578_p2 = (tmp_202_fu_9518_p3 ^ tmp_200_fu_9496_p3);

assign xor_ln65_8_fu_9584_p2 = (xor_ln65_7_fu_9578_p2 ^ xor_ln65_6_fu_9572_p2);

assign xor_ln65_9_fu_9714_p2 = (tmp_212_fu_9706_p3 ^ tmp_211_fu_9698_p3);

assign xor_ln65_fu_3236_p2 = (tmp_67_fu_3228_p3 ^ tmp_66_fu_3220_p3);

assign xor_ln70_fu_9756_p2 = (res_39_fu_9742_p6 ^ a0_fu_9604_p2);

assign xor_ln86_10_fu_1304_p2 = (and_ln86_15_fu_1292_p2 ^ and_ln86_14_fu_1270_p2);

assign xor_ln86_11_fu_1310_p2 = (xor_ln86_9_fu_1298_p2 ^ xor_ln86_10_fu_1304_p2);

assign xor_ln86_12_fu_1612_p2 = (and_ln86_17_fu_1562_p2 ^ and_ln86_16_fu_1540_p2);

assign xor_ln86_13_fu_1618_p2 = (and_ln86_19_fu_1606_p2 ^ and_ln86_18_fu_1584_p2);

assign xor_ln86_14_fu_1624_p2 = (xor_ln86_13_fu_1618_p2 ^ xor_ln86_12_fu_1612_p2);

assign xor_ln86_15_fu_1910_p2 = (and_ln86_22_fu_1882_p2 ^ and_ln86_21_fu_1860_p2);

assign xor_ln86_16_fu_1916_p2 = (and_ln86_23_fu_1904_p2 ^ and_ln86_20_fu_1838_p2);

assign xor_ln86_17_fu_1922_p2 = (xor_ln86_16_fu_1916_p2 ^ xor_ln86_15_fu_1910_p2);

assign xor_ln86_18_fu_2290_p2 = (and_ln86_25_fu_2240_p2 ^ and_ln86_24_fu_2218_p2);

assign xor_ln86_19_fu_2296_p2 = (and_ln86_27_fu_2284_p2 ^ and_ln86_26_fu_2262_p2);

assign xor_ln86_1_fu_300_p2 = (and_ln86_3_fu_288_p2 ^ and_ln86_2_fu_266_p2);

assign xor_ln86_20_fu_2302_p2 = (xor_ln86_19_fu_2296_p2 ^ xor_ln86_18_fu_2290_p2);

assign xor_ln86_21_fu_2592_p2 = (and_ln86_29_fu_2542_p2 ^ and_ln86_28_fu_2520_p2);

assign xor_ln86_22_fu_2598_p2 = (and_ln86_31_fu_2586_p2 ^ and_ln86_30_fu_2564_p2);

assign xor_ln86_23_fu_2604_p2 = (xor_ln86_22_fu_2598_p2 ^ xor_ln86_21_fu_2592_p2);

assign xor_ln86_24_fu_2890_p2 = (and_ln86_34_fu_2862_p2 ^ and_ln86_33_fu_2840_p2);

assign xor_ln86_25_fu_2896_p2 = (and_ln86_35_fu_2884_p2 ^ and_ln86_32_fu_2818_p2);

assign xor_ln86_26_fu_2902_p2 = (xor_ln86_25_fu_2896_p2 ^ xor_ln86_24_fu_2890_p2);

assign xor_ln86_27_fu_3496_p2 = (and_ln86_37_fu_3446_p2 ^ and_ln86_36_fu_3424_p2);

assign xor_ln86_28_fu_3502_p2 = (and_ln86_39_fu_3490_p2 ^ and_ln86_38_fu_3468_p2);

assign xor_ln86_29_fu_3508_p2 = (xor_ln86_28_fu_3502_p2 ^ xor_ln86_27_fu_3496_p2);

assign xor_ln86_2_fu_306_p2 = (xor_ln86_fu_294_p2 ^ xor_ln86_1_fu_300_p2);

assign xor_ln86_30_fu_3798_p2 = (and_ln86_41_fu_3748_p2 ^ and_ln86_40_fu_3726_p2);

assign xor_ln86_31_fu_3804_p2 = (and_ln86_43_fu_3792_p2 ^ and_ln86_42_fu_3770_p2);

assign xor_ln86_32_fu_3810_p2 = (xor_ln86_31_fu_3804_p2 ^ xor_ln86_30_fu_3798_p2);

assign xor_ln86_33_fu_4096_p2 = (and_ln86_46_fu_4068_p2 ^ and_ln86_45_fu_4046_p2);

assign xor_ln86_34_fu_4102_p2 = (and_ln86_47_fu_4090_p2 ^ and_ln86_44_fu_4024_p2);

assign xor_ln86_35_fu_4108_p2 = (xor_ln86_34_fu_4102_p2 ^ xor_ln86_33_fu_4096_p2);

assign xor_ln86_36_fu_4500_p2 = (and_ln86_49_fu_4450_p2 ^ and_ln86_48_fu_4428_p2);

assign xor_ln86_37_fu_4506_p2 = (and_ln86_51_fu_4494_p2 ^ and_ln86_50_fu_4472_p2);

assign xor_ln86_38_fu_4512_p2 = (xor_ln86_37_fu_4506_p2 ^ xor_ln86_36_fu_4500_p2);

assign xor_ln86_39_fu_4814_p2 = (and_ln86_53_fu_4764_p2 ^ and_ln86_52_fu_4742_p2);

assign xor_ln86_3_fu_596_p2 = (and_ln86_5_fu_546_p2 ^ and_ln86_4_fu_524_p2);

assign xor_ln86_40_fu_4820_p2 = (and_ln86_55_fu_4808_p2 ^ and_ln86_54_fu_4786_p2);

assign xor_ln86_41_fu_4826_p2 = (xor_ln86_40_fu_4820_p2 ^ xor_ln86_39_fu_4814_p2);

assign xor_ln86_42_fu_5112_p2 = (and_ln86_58_fu_5084_p2 ^ and_ln86_57_fu_5062_p2);

assign xor_ln86_43_fu_5118_p2 = (and_ln86_59_fu_5106_p2 ^ and_ln86_56_fu_5040_p2);

assign xor_ln86_44_fu_5124_p2 = (xor_ln86_43_fu_5118_p2 ^ xor_ln86_42_fu_5112_p2);

assign xor_ln86_45_fu_5492_p2 = (and_ln86_61_fu_5442_p2 ^ and_ln86_60_fu_5420_p2);

assign xor_ln86_46_fu_5498_p2 = (and_ln86_63_fu_5486_p2 ^ and_ln86_62_fu_5464_p2);

assign xor_ln86_47_fu_5504_p2 = (xor_ln86_46_fu_5498_p2 ^ xor_ln86_45_fu_5492_p2);

assign xor_ln86_48_fu_5794_p2 = (and_ln86_65_fu_5744_p2 ^ and_ln86_64_fu_5722_p2);

assign xor_ln86_49_fu_5800_p2 = (and_ln86_67_fu_5788_p2 ^ and_ln86_66_fu_5766_p2);

assign xor_ln86_4_fu_602_p2 = (and_ln86_7_fu_590_p2 ^ and_ln86_6_fu_568_p2);

assign xor_ln86_50_fu_5806_p2 = (xor_ln86_49_fu_5800_p2 ^ xor_ln86_48_fu_5794_p2);

assign xor_ln86_51_fu_6092_p2 = (and_ln86_70_fu_6064_p2 ^ and_ln86_69_fu_6042_p2);

assign xor_ln86_52_fu_6098_p2 = (and_ln86_71_fu_6086_p2 ^ and_ln86_68_fu_6020_p2);

assign xor_ln86_53_fu_6104_p2 = (xor_ln86_52_fu_6098_p2 ^ xor_ln86_51_fu_6092_p2);

assign xor_ln86_54_fu_6630_p2 = (and_ln86_73_fu_6580_p2 ^ and_ln86_72_fu_6558_p2);

assign xor_ln86_55_fu_6636_p2 = (and_ln86_75_fu_6624_p2 ^ and_ln86_74_fu_6602_p2);

assign xor_ln86_56_fu_6642_p2 = (xor_ln86_55_fu_6636_p2 ^ xor_ln86_54_fu_6630_p2);

assign xor_ln86_57_fu_6932_p2 = (and_ln86_77_fu_6882_p2 ^ and_ln86_76_fu_6860_p2);

assign xor_ln86_58_fu_6938_p2 = (and_ln86_79_fu_6926_p2 ^ and_ln86_78_fu_6904_p2);

assign xor_ln86_59_fu_6944_p2 = (xor_ln86_58_fu_6938_p2 ^ xor_ln86_57_fu_6932_p2);

assign xor_ln86_5_fu_608_p2 = (xor_ln86_4_fu_602_p2 ^ xor_ln86_3_fu_596_p2);

assign xor_ln86_60_fu_7230_p2 = (and_ln86_82_fu_7202_p2 ^ and_ln86_81_fu_7180_p2);

assign xor_ln86_61_fu_7236_p2 = (and_ln86_83_fu_7224_p2 ^ and_ln86_80_fu_7158_p2);

assign xor_ln86_62_fu_7242_p2 = (xor_ln86_61_fu_7236_p2 ^ xor_ln86_60_fu_7230_p2);

assign xor_ln86_63_fu_7634_p2 = (and_ln86_85_fu_7584_p2 ^ and_ln86_84_fu_7562_p2);

assign xor_ln86_64_fu_7640_p2 = (and_ln86_87_fu_7628_p2 ^ and_ln86_86_fu_7606_p2);

assign xor_ln86_65_fu_7646_p2 = (xor_ln86_64_fu_7640_p2 ^ xor_ln86_63_fu_7634_p2);

assign xor_ln86_66_fu_7948_p2 = (and_ln86_89_fu_7898_p2 ^ and_ln86_88_fu_7876_p2);

assign xor_ln86_67_fu_7954_p2 = (and_ln86_91_fu_7942_p2 ^ and_ln86_90_fu_7920_p2);

assign xor_ln86_68_fu_7960_p2 = (xor_ln86_67_fu_7954_p2 ^ xor_ln86_66_fu_7948_p2);

assign xor_ln86_69_fu_8246_p2 = (and_ln86_94_fu_8218_p2 ^ and_ln86_93_fu_8196_p2);

assign xor_ln86_6_fu_894_p2 = (and_ln86_9_fu_844_p2 ^ and_ln86_10_fu_866_p2);

assign xor_ln86_70_fu_8252_p2 = (and_ln86_95_fu_8240_p2 ^ and_ln86_92_fu_8174_p2);

assign xor_ln86_71_fu_8258_p2 = (xor_ln86_70_fu_8252_p2 ^ xor_ln86_69_fu_8246_p2);

assign xor_ln86_72_fu_8626_p2 = (and_ln86_97_fu_8576_p2 ^ and_ln86_96_fu_8554_p2);

assign xor_ln86_73_fu_8632_p2 = (and_ln86_99_fu_8620_p2 ^ and_ln86_98_fu_8598_p2);

assign xor_ln86_74_fu_8638_p2 = (xor_ln86_73_fu_8632_p2 ^ xor_ln86_72_fu_8626_p2);

assign xor_ln86_75_fu_8928_p2 = (and_ln86_101_fu_8878_p2 ^ and_ln86_100_fu_8856_p2);

assign xor_ln86_76_fu_8934_p2 = (and_ln86_103_fu_8922_p2 ^ and_ln86_102_fu_8900_p2);

assign xor_ln86_77_fu_8940_p2 = (xor_ln86_76_fu_8934_p2 ^ xor_ln86_75_fu_8928_p2);

assign xor_ln86_78_fu_9226_p2 = (and_ln86_106_fu_9198_p2 ^ and_ln86_105_fu_9176_p2);

assign xor_ln86_79_fu_9232_p2 = (and_ln86_107_fu_9220_p2 ^ and_ln86_104_fu_9154_p2);

assign xor_ln86_7_fu_900_p2 = (and_ln86_8_fu_822_p2 ^ and_ln86_11_fu_888_p2);

assign xor_ln86_80_fu_9238_p2 = (xor_ln86_79_fu_9232_p2 ^ xor_ln86_78_fu_9226_p2);

assign xor_ln86_8_fu_906_p2 = (xor_ln86_7_fu_900_p2 ^ xor_ln86_6_fu_894_p2);

assign xor_ln86_9_fu_1298_p2 = (and_ln86_13_fu_1248_p2 ^ and_ln86_12_fu_1226_p2);

assign xor_ln86_fu_294_p2 = (and_ln86_fu_222_p2 ^ and_ln86_1_fu_244_p2);

assign xor_ln87_100_fu_7266_p2 = (and_ln87_81_fu_7254_p2 ^ and_ln86_81_fu_7180_p2);

assign xor_ln87_101_fu_7272_p2 = (and_ln87_82_fu_7260_p2 ^ and_ln87_80_fu_7248_p2);

assign xor_ln87_102_fu_7278_p2 = (xor_ln87_101_fu_7272_p2 ^ xor_ln87_100_fu_7266_p2);

assign xor_ln87_103_fu_7290_p2 = (and_ln87_83_fu_7284_p2 ^ and_ln86_83_fu_7224_p2);

assign xor_ln87_104_fu_7296_p2 = (xor_ln87_103_fu_7290_p2 ^ xor_ln87_102_fu_7278_p2);

assign xor_ln87_105_fu_7676_p2 = (and_ln87_85_fu_7658_p2 ^ and_ln86_85_fu_7584_p2);

assign xor_ln87_106_fu_7682_p2 = (xor_ln87_105_fu_7676_p2 ^ and_ln87_84_fu_7652_p2);

assign xor_ln87_107_fu_7688_p2 = (and_ln87_87_fu_7670_p2 ^ and_ln86_87_fu_7628_p2);

assign xor_ln87_108_fu_7694_p2 = (xor_ln87_107_fu_7688_p2 ^ and_ln87_86_fu_7664_p2);

assign xor_ln87_109_fu_7700_p2 = (xor_ln87_108_fu_7694_p2 ^ xor_ln87_106_fu_7682_p2);

assign xor_ln87_10_fu_930_p2 = (and_ln87_9_fu_918_p2 ^ and_ln86_9_fu_844_p2);

assign xor_ln87_110_fu_7990_p2 = (and_ln87_89_fu_7972_p2 ^ and_ln86_89_fu_7898_p2);

assign xor_ln87_111_fu_7996_p2 = (xor_ln87_110_fu_7990_p2 ^ and_ln87_88_fu_7966_p2);

assign xor_ln87_112_fu_8002_p2 = (and_ln87_91_fu_7984_p2 ^ and_ln86_91_fu_7942_p2);

assign xor_ln87_113_fu_8008_p2 = (xor_ln87_112_fu_8002_p2 ^ and_ln87_90_fu_7978_p2);

assign xor_ln87_114_fu_8014_p2 = (xor_ln87_113_fu_8008_p2 ^ xor_ln87_111_fu_7996_p2);

assign xor_ln87_115_fu_8282_p2 = (and_ln87_93_fu_8270_p2 ^ and_ln86_93_fu_8196_p2);

assign xor_ln87_116_fu_8288_p2 = (and_ln87_94_fu_8276_p2 ^ and_ln87_92_fu_8264_p2);

assign xor_ln87_117_fu_8294_p2 = (xor_ln87_116_fu_8288_p2 ^ xor_ln87_115_fu_8282_p2);

assign xor_ln87_118_fu_8306_p2 = (and_ln87_95_fu_8300_p2 ^ and_ln86_95_fu_8240_p2);

assign xor_ln87_119_fu_8312_p2 = (xor_ln87_118_fu_8306_p2 ^ xor_ln87_117_fu_8294_p2);

assign xor_ln87_11_fu_936_p2 = (and_ln87_8_fu_912_p2 ^ and_ln87_10_fu_924_p2);

assign xor_ln87_120_fu_8668_p2 = (and_ln87_97_fu_8650_p2 ^ and_ln86_97_fu_8576_p2);

assign xor_ln87_121_fu_8674_p2 = (xor_ln87_120_fu_8668_p2 ^ and_ln87_96_fu_8644_p2);

assign xor_ln87_122_fu_8680_p2 = (and_ln87_99_fu_8662_p2 ^ and_ln86_99_fu_8620_p2);

assign xor_ln87_123_fu_8686_p2 = (xor_ln87_122_fu_8680_p2 ^ and_ln87_98_fu_8656_p2);

assign xor_ln87_124_fu_8692_p2 = (xor_ln87_123_fu_8686_p2 ^ xor_ln87_121_fu_8674_p2);

assign xor_ln87_125_fu_8970_p2 = (and_ln87_101_fu_8952_p2 ^ and_ln86_101_fu_8878_p2);

assign xor_ln87_126_fu_8976_p2 = (xor_ln87_125_fu_8970_p2 ^ and_ln87_100_fu_8946_p2);

assign xor_ln87_127_fu_8982_p2 = (and_ln87_103_fu_8964_p2 ^ and_ln86_103_fu_8922_p2);

assign xor_ln87_128_fu_8988_p2 = (xor_ln87_127_fu_8982_p2 ^ and_ln87_102_fu_8958_p2);

assign xor_ln87_129_fu_8994_p2 = (xor_ln87_128_fu_8988_p2 ^ xor_ln87_126_fu_8976_p2);

assign xor_ln87_12_fu_942_p2 = (xor_ln87_11_fu_936_p2 ^ xor_ln87_10_fu_930_p2);

assign xor_ln87_130_fu_9262_p2 = (and_ln87_105_fu_9250_p2 ^ and_ln86_105_fu_9176_p2);

assign xor_ln87_131_fu_9268_p2 = (and_ln87_106_fu_9256_p2 ^ and_ln87_104_fu_9244_p2);

assign xor_ln87_132_fu_9274_p2 = (xor_ln87_131_fu_9268_p2 ^ xor_ln87_130_fu_9262_p2);

assign xor_ln87_133_fu_9286_p2 = (and_ln87_107_fu_9280_p2 ^ and_ln86_107_fu_9220_p2);

assign xor_ln87_134_fu_9292_p2 = (xor_ln87_133_fu_9286_p2 ^ xor_ln87_132_fu_9274_p2);

assign xor_ln87_13_fu_954_p2 = (and_ln87_11_fu_948_p2 ^ and_ln86_11_fu_888_p2);

assign xor_ln87_14_fu_960_p2 = (xor_ln87_13_fu_954_p2 ^ xor_ln87_12_fu_942_p2);

assign xor_ln87_15_fu_1340_p2 = (and_ln87_13_fu_1322_p2 ^ and_ln86_13_fu_1248_p2);

assign xor_ln87_16_fu_1346_p2 = (xor_ln87_15_fu_1340_p2 ^ and_ln87_12_fu_1316_p2);

assign xor_ln87_17_fu_1352_p2 = (and_ln87_15_fu_1334_p2 ^ and_ln86_15_fu_1292_p2);

assign xor_ln87_18_fu_1358_p2 = (xor_ln87_17_fu_1352_p2 ^ and_ln87_14_fu_1328_p2);

assign xor_ln87_19_fu_1364_p2 = (xor_ln87_18_fu_1358_p2 ^ xor_ln87_16_fu_1346_p2);

assign xor_ln87_1_fu_342_p2 = (xor_ln87_fu_336_p2 ^ and_ln87_fu_312_p2);

assign xor_ln87_20_fu_1654_p2 = (and_ln87_17_fu_1636_p2 ^ and_ln86_17_fu_1562_p2);

assign xor_ln87_21_fu_1660_p2 = (xor_ln87_20_fu_1654_p2 ^ and_ln87_16_fu_1630_p2);

assign xor_ln87_22_fu_1666_p2 = (and_ln87_19_fu_1648_p2 ^ and_ln86_19_fu_1606_p2);

assign xor_ln87_23_fu_1672_p2 = (xor_ln87_22_fu_1666_p2 ^ and_ln87_18_fu_1642_p2);

assign xor_ln87_24_fu_1678_p2 = (xor_ln87_23_fu_1672_p2 ^ xor_ln87_21_fu_1660_p2);

assign xor_ln87_25_fu_1946_p2 = (and_ln87_21_fu_1934_p2 ^ and_ln86_21_fu_1860_p2);

assign xor_ln87_26_fu_1952_p2 = (and_ln87_22_fu_1940_p2 ^ and_ln87_20_fu_1928_p2);

assign xor_ln87_27_fu_1958_p2 = (xor_ln87_26_fu_1952_p2 ^ xor_ln87_25_fu_1946_p2);

assign xor_ln87_28_fu_1970_p2 = (and_ln87_23_fu_1964_p2 ^ and_ln86_23_fu_1904_p2);

assign xor_ln87_29_fu_1976_p2 = (xor_ln87_28_fu_1970_p2 ^ xor_ln87_27_fu_1958_p2);

assign xor_ln87_2_fu_348_p2 = (and_ln87_3_fu_330_p2 ^ and_ln86_3_fu_288_p2);

assign xor_ln87_30_fu_2332_p2 = (and_ln87_25_fu_2314_p2 ^ and_ln86_25_fu_2240_p2);

assign xor_ln87_31_fu_2338_p2 = (xor_ln87_30_fu_2332_p2 ^ and_ln87_24_fu_2308_p2);

assign xor_ln87_32_fu_2344_p2 = (and_ln87_27_fu_2326_p2 ^ and_ln86_27_fu_2284_p2);

assign xor_ln87_33_fu_2350_p2 = (xor_ln87_32_fu_2344_p2 ^ and_ln87_26_fu_2320_p2);

assign xor_ln87_34_fu_2356_p2 = (xor_ln87_33_fu_2350_p2 ^ xor_ln87_31_fu_2338_p2);

assign xor_ln87_35_fu_2634_p2 = (and_ln87_29_fu_2616_p2 ^ and_ln86_29_fu_2542_p2);

assign xor_ln87_36_fu_2640_p2 = (xor_ln87_35_fu_2634_p2 ^ and_ln87_28_fu_2610_p2);

assign xor_ln87_37_fu_2646_p2 = (and_ln87_31_fu_2628_p2 ^ and_ln86_31_fu_2586_p2);

assign xor_ln87_38_fu_2652_p2 = (xor_ln87_37_fu_2646_p2 ^ and_ln87_30_fu_2622_p2);

assign xor_ln87_39_fu_2658_p2 = (xor_ln87_38_fu_2652_p2 ^ xor_ln87_36_fu_2640_p2);

assign xor_ln87_3_fu_354_p2 = (xor_ln87_2_fu_348_p2 ^ and_ln87_2_fu_324_p2);

assign xor_ln87_40_fu_2926_p2 = (and_ln87_33_fu_2914_p2 ^ and_ln86_33_fu_2840_p2);

assign xor_ln87_41_fu_2932_p2 = (and_ln87_34_fu_2920_p2 ^ and_ln87_32_fu_2908_p2);

assign xor_ln87_42_fu_2938_p2 = (xor_ln87_41_fu_2932_p2 ^ xor_ln87_40_fu_2926_p2);

assign xor_ln87_43_fu_2950_p2 = (and_ln87_35_fu_2944_p2 ^ and_ln86_35_fu_2884_p2);

assign xor_ln87_44_fu_2956_p2 = (xor_ln87_43_fu_2950_p2 ^ xor_ln87_42_fu_2938_p2);

assign xor_ln87_45_fu_3538_p2 = (and_ln87_37_fu_3520_p2 ^ and_ln86_37_fu_3446_p2);

assign xor_ln87_46_fu_3544_p2 = (xor_ln87_45_fu_3538_p2 ^ and_ln87_36_fu_3514_p2);

assign xor_ln87_47_fu_3550_p2 = (and_ln87_39_fu_3532_p2 ^ and_ln86_39_fu_3490_p2);

assign xor_ln87_48_fu_3556_p2 = (xor_ln87_47_fu_3550_p2 ^ and_ln87_38_fu_3526_p2);

assign xor_ln87_49_fu_3562_p2 = (xor_ln87_48_fu_3556_p2 ^ xor_ln87_46_fu_3544_p2);

assign xor_ln87_4_fu_360_p2 = (xor_ln87_3_fu_354_p2 ^ xor_ln87_1_fu_342_p2);

assign xor_ln87_50_fu_3840_p2 = (and_ln87_41_fu_3822_p2 ^ and_ln86_41_fu_3748_p2);

assign xor_ln87_51_fu_3846_p2 = (xor_ln87_50_fu_3840_p2 ^ and_ln87_40_fu_3816_p2);

assign xor_ln87_52_fu_3852_p2 = (and_ln87_43_fu_3834_p2 ^ and_ln86_43_fu_3792_p2);

assign xor_ln87_53_fu_3858_p2 = (xor_ln87_52_fu_3852_p2 ^ and_ln87_42_fu_3828_p2);

assign xor_ln87_54_fu_3864_p2 = (xor_ln87_53_fu_3858_p2 ^ xor_ln87_51_fu_3846_p2);

assign xor_ln87_55_fu_4132_p2 = (and_ln87_45_fu_4120_p2 ^ and_ln86_45_fu_4046_p2);

assign xor_ln87_56_fu_4138_p2 = (and_ln87_46_fu_4126_p2 ^ and_ln87_44_fu_4114_p2);

assign xor_ln87_57_fu_4144_p2 = (xor_ln87_56_fu_4138_p2 ^ xor_ln87_55_fu_4132_p2);

assign xor_ln87_58_fu_4156_p2 = (and_ln87_47_fu_4150_p2 ^ and_ln86_47_fu_4090_p2);

assign xor_ln87_59_fu_4162_p2 = (xor_ln87_58_fu_4156_p2 ^ xor_ln87_57_fu_4144_p2);

assign xor_ln87_5_fu_638_p2 = (and_ln87_5_fu_620_p2 ^ and_ln86_5_fu_546_p2);

assign xor_ln87_60_fu_4542_p2 = (and_ln87_49_fu_4524_p2 ^ and_ln86_49_fu_4450_p2);

assign xor_ln87_61_fu_4548_p2 = (xor_ln87_60_fu_4542_p2 ^ and_ln87_48_fu_4518_p2);

assign xor_ln87_62_fu_4554_p2 = (and_ln87_51_fu_4536_p2 ^ and_ln86_51_fu_4494_p2);

assign xor_ln87_63_fu_4560_p2 = (xor_ln87_62_fu_4554_p2 ^ and_ln87_50_fu_4530_p2);

assign xor_ln87_64_fu_4566_p2 = (xor_ln87_63_fu_4560_p2 ^ xor_ln87_61_fu_4548_p2);

assign xor_ln87_65_fu_4856_p2 = (and_ln87_53_fu_4838_p2 ^ and_ln86_53_fu_4764_p2);

assign xor_ln87_66_fu_4862_p2 = (xor_ln87_65_fu_4856_p2 ^ and_ln87_52_fu_4832_p2);

assign xor_ln87_67_fu_4868_p2 = (and_ln87_55_fu_4850_p2 ^ and_ln86_55_fu_4808_p2);

assign xor_ln87_68_fu_4874_p2 = (xor_ln87_67_fu_4868_p2 ^ and_ln87_54_fu_4844_p2);

assign xor_ln87_69_fu_4880_p2 = (xor_ln87_68_fu_4874_p2 ^ xor_ln87_66_fu_4862_p2);

assign xor_ln87_6_fu_644_p2 = (xor_ln87_5_fu_638_p2 ^ and_ln87_4_fu_614_p2);

assign xor_ln87_70_fu_5148_p2 = (and_ln87_57_fu_5136_p2 ^ and_ln86_57_fu_5062_p2);

assign xor_ln87_71_fu_5154_p2 = (and_ln87_58_fu_5142_p2 ^ and_ln87_56_fu_5130_p2);

assign xor_ln87_72_fu_5160_p2 = (xor_ln87_71_fu_5154_p2 ^ xor_ln87_70_fu_5148_p2);

assign xor_ln87_73_fu_5172_p2 = (and_ln87_59_fu_5166_p2 ^ and_ln86_59_fu_5106_p2);

assign xor_ln87_74_fu_5178_p2 = (xor_ln87_73_fu_5172_p2 ^ xor_ln87_72_fu_5160_p2);

assign xor_ln87_75_fu_5534_p2 = (and_ln87_61_fu_5516_p2 ^ and_ln86_61_fu_5442_p2);

assign xor_ln87_76_fu_5540_p2 = (xor_ln87_75_fu_5534_p2 ^ and_ln87_60_fu_5510_p2);

assign xor_ln87_77_fu_5546_p2 = (and_ln87_63_fu_5528_p2 ^ and_ln86_63_fu_5486_p2);

assign xor_ln87_78_fu_5552_p2 = (xor_ln87_77_fu_5546_p2 ^ and_ln87_62_fu_5522_p2);

assign xor_ln87_79_fu_5558_p2 = (xor_ln87_78_fu_5552_p2 ^ xor_ln87_76_fu_5540_p2);

assign xor_ln87_7_fu_650_p2 = (and_ln87_7_fu_632_p2 ^ and_ln86_7_fu_590_p2);

assign xor_ln87_80_fu_5836_p2 = (and_ln87_65_fu_5818_p2 ^ and_ln86_65_fu_5744_p2);

assign xor_ln87_81_fu_5842_p2 = (xor_ln87_80_fu_5836_p2 ^ and_ln87_64_fu_5812_p2);

assign xor_ln87_82_fu_5848_p2 = (and_ln87_67_fu_5830_p2 ^ and_ln86_67_fu_5788_p2);

assign xor_ln87_83_fu_5854_p2 = (xor_ln87_82_fu_5848_p2 ^ and_ln87_66_fu_5824_p2);

assign xor_ln87_84_fu_5860_p2 = (xor_ln87_83_fu_5854_p2 ^ xor_ln87_81_fu_5842_p2);

assign xor_ln87_85_fu_6128_p2 = (and_ln87_69_fu_6116_p2 ^ and_ln86_69_fu_6042_p2);

assign xor_ln87_86_fu_6134_p2 = (and_ln87_70_fu_6122_p2 ^ and_ln87_68_fu_6110_p2);

assign xor_ln87_87_fu_6140_p2 = (xor_ln87_86_fu_6134_p2 ^ xor_ln87_85_fu_6128_p2);

assign xor_ln87_88_fu_6152_p2 = (and_ln87_71_fu_6146_p2 ^ and_ln86_71_fu_6086_p2);

assign xor_ln87_89_fu_6158_p2 = (xor_ln87_88_fu_6152_p2 ^ xor_ln87_87_fu_6140_p2);

assign xor_ln87_8_fu_656_p2 = (xor_ln87_7_fu_650_p2 ^ and_ln87_6_fu_626_p2);

assign xor_ln87_90_fu_6672_p2 = (and_ln87_73_fu_6654_p2 ^ and_ln86_73_fu_6580_p2);

assign xor_ln87_91_fu_6678_p2 = (xor_ln87_90_fu_6672_p2 ^ and_ln87_72_fu_6648_p2);

assign xor_ln87_92_fu_6684_p2 = (and_ln87_75_fu_6666_p2 ^ and_ln86_75_fu_6624_p2);

assign xor_ln87_93_fu_6690_p2 = (xor_ln87_92_fu_6684_p2 ^ and_ln87_74_fu_6660_p2);

assign xor_ln87_94_fu_6696_p2 = (xor_ln87_93_fu_6690_p2 ^ xor_ln87_91_fu_6678_p2);

assign xor_ln87_95_fu_6974_p2 = (and_ln87_77_fu_6956_p2 ^ and_ln86_77_fu_6882_p2);

assign xor_ln87_96_fu_6980_p2 = (xor_ln87_95_fu_6974_p2 ^ and_ln87_76_fu_6950_p2);

assign xor_ln87_97_fu_6986_p2 = (and_ln87_79_fu_6968_p2 ^ and_ln86_79_fu_6926_p2);

assign xor_ln87_98_fu_6992_p2 = (xor_ln87_97_fu_6986_p2 ^ and_ln87_78_fu_6962_p2);

assign xor_ln87_99_fu_6998_p2 = (xor_ln87_98_fu_6992_p2 ^ xor_ln87_96_fu_6980_p2);

assign xor_ln87_9_fu_662_p2 = (xor_ln87_8_fu_656_p2 ^ xor_ln87_6_fu_644_p2);

assign xor_ln87_fu_336_p2 = (and_ln87_1_fu_318_p2 ^ and_ln86_1_fu_244_p2);

assign xor_ln88_100_fu_7326_p2 = (and_ln88_82_fu_7314_p2 ^ and_ln87_82_fu_7260_p2);

assign xor_ln88_101_fu_7332_p2 = (and_ln88_83_fu_7320_p2 ^ and_ln88_80_fu_7302_p2);

assign xor_ln88_102_fu_7338_p2 = (xor_ln88_101_fu_7332_p2 ^ and_ln88_81_fu_7308_p2);

assign xor_ln88_103_fu_7344_p2 = (xor_ln88_102_fu_7338_p2 ^ xor_ln88_100_fu_7326_p2);

assign xor_ln88_104_fu_7350_p2 = (xor_ln88_103_fu_7344_p2 ^ xor_ln87_103_fu_7290_p2);

assign xor_ln88_105_fu_7730_p2 = (and_ln88_86_fu_7718_p2 ^ and_ln88_85_fu_7712_p2);

assign xor_ln88_106_fu_7736_p2 = (xor_ln88_105_fu_7730_p2 ^ and_ln88_84_fu_7706_p2);

assign xor_ln88_107_fu_7742_p2 = (and_ln88_87_fu_7724_p2 ^ and_ln87_86_fu_7664_p2);

assign xor_ln88_108_fu_7748_p2 = (xor_ln88_107_fu_7742_p2 ^ xor_ln87_107_fu_7688_p2);

assign xor_ln88_109_fu_7754_p2 = (xor_ln88_108_fu_7748_p2 ^ xor_ln88_106_fu_7736_p2);

assign xor_ln88_10_fu_990_p2 = (and_ln88_10_fu_978_p2 ^ and_ln87_10_fu_924_p2);

assign xor_ln88_110_fu_8044_p2 = (and_ln88_90_fu_8032_p2 ^ and_ln88_89_fu_8026_p2);

assign xor_ln88_111_fu_8050_p2 = (xor_ln88_110_fu_8044_p2 ^ and_ln88_88_fu_8020_p2);

assign xor_ln88_112_fu_8056_p2 = (and_ln88_91_fu_8038_p2 ^ and_ln87_90_fu_7978_p2);

assign xor_ln88_113_fu_8062_p2 = (xor_ln88_112_fu_8056_p2 ^ xor_ln87_112_fu_8002_p2);

assign xor_ln88_114_fu_8068_p2 = (xor_ln88_113_fu_8062_p2 ^ xor_ln88_111_fu_8050_p2);

assign xor_ln88_115_fu_8342_p2 = (and_ln88_94_fu_8330_p2 ^ and_ln87_94_fu_8276_p2);

assign xor_ln88_116_fu_8348_p2 = (and_ln88_95_fu_8336_p2 ^ and_ln88_92_fu_8318_p2);

assign xor_ln88_117_fu_8354_p2 = (xor_ln88_116_fu_8348_p2 ^ and_ln88_93_fu_8324_p2);

assign xor_ln88_118_fu_8360_p2 = (xor_ln88_117_fu_8354_p2 ^ xor_ln88_115_fu_8342_p2);

assign xor_ln88_119_fu_8366_p2 = (xor_ln88_118_fu_8360_p2 ^ xor_ln87_118_fu_8306_p2);

assign xor_ln88_11_fu_996_p2 = (and_ln88_8_fu_966_p2 ^ and_ln88_11_fu_984_p2);

assign xor_ln88_120_fu_8722_p2 = (and_ln88_98_fu_8710_p2 ^ and_ln88_97_fu_8704_p2);

assign xor_ln88_121_fu_8728_p2 = (xor_ln88_120_fu_8722_p2 ^ and_ln88_96_fu_8698_p2);

assign xor_ln88_122_fu_8734_p2 = (and_ln88_99_fu_8716_p2 ^ and_ln87_98_fu_8656_p2);

assign xor_ln88_123_fu_8740_p2 = (xor_ln88_122_fu_8734_p2 ^ xor_ln87_122_fu_8680_p2);

assign xor_ln88_124_fu_8746_p2 = (xor_ln88_123_fu_8740_p2 ^ xor_ln88_121_fu_8728_p2);

assign xor_ln88_125_fu_9024_p2 = (and_ln88_102_fu_9012_p2 ^ and_ln88_101_fu_9006_p2);

assign xor_ln88_126_fu_9030_p2 = (xor_ln88_125_fu_9024_p2 ^ and_ln88_100_fu_9000_p2);

assign xor_ln88_127_fu_9036_p2 = (and_ln88_103_fu_9018_p2 ^ and_ln87_102_fu_8958_p2);

assign xor_ln88_128_fu_9042_p2 = (xor_ln88_127_fu_9036_p2 ^ xor_ln87_127_fu_8982_p2);

assign xor_ln88_129_fu_9048_p2 = (xor_ln88_128_fu_9042_p2 ^ xor_ln88_126_fu_9030_p2);

assign xor_ln88_12_fu_1002_p2 = (xor_ln88_11_fu_996_p2 ^ and_ln88_9_fu_972_p2);

assign xor_ln88_130_fu_9322_p2 = (and_ln88_106_fu_9310_p2 ^ and_ln87_106_fu_9256_p2);

assign xor_ln88_131_fu_9328_p2 = (and_ln88_107_fu_9316_p2 ^ and_ln88_104_fu_9298_p2);

assign xor_ln88_132_fu_9334_p2 = (xor_ln88_131_fu_9328_p2 ^ and_ln88_105_fu_9304_p2);

assign xor_ln88_133_fu_9340_p2 = (xor_ln88_132_fu_9334_p2 ^ xor_ln88_130_fu_9322_p2);

assign xor_ln88_134_fu_9346_p2 = (xor_ln88_133_fu_9340_p2 ^ xor_ln87_133_fu_9286_p2);

assign xor_ln88_13_fu_1008_p2 = (xor_ln88_12_fu_1002_p2 ^ xor_ln88_10_fu_990_p2);

assign xor_ln88_14_fu_1014_p2 = (xor_ln88_13_fu_1008_p2 ^ xor_ln87_13_fu_954_p2);

assign xor_ln88_15_fu_1394_p2 = (and_ln88_14_fu_1382_p2 ^ and_ln88_13_fu_1376_p2);

assign xor_ln88_16_fu_1400_p2 = (xor_ln88_15_fu_1394_p2 ^ and_ln88_12_fu_1370_p2);

assign xor_ln88_17_fu_1406_p2 = (and_ln88_15_fu_1388_p2 ^ and_ln87_14_fu_1328_p2);

assign xor_ln88_18_fu_1412_p2 = (xor_ln88_17_fu_1406_p2 ^ xor_ln87_17_fu_1352_p2);

assign xor_ln88_19_fu_1418_p2 = (xor_ln88_18_fu_1412_p2 ^ xor_ln88_16_fu_1400_p2);

assign xor_ln88_1_fu_396_p2 = (xor_ln88_fu_390_p2 ^ and_ln88_fu_366_p2);

assign xor_ln88_20_fu_1708_p2 = (and_ln88_18_fu_1696_p2 ^ and_ln88_17_fu_1690_p2);

assign xor_ln88_21_fu_1714_p2 = (xor_ln88_20_fu_1708_p2 ^ and_ln88_16_fu_1684_p2);

assign xor_ln88_22_fu_1720_p2 = (and_ln88_19_fu_1702_p2 ^ and_ln87_18_fu_1642_p2);

assign xor_ln88_23_fu_1726_p2 = (xor_ln88_22_fu_1720_p2 ^ xor_ln87_22_fu_1666_p2);

assign xor_ln88_24_fu_1732_p2 = (xor_ln88_23_fu_1726_p2 ^ xor_ln88_21_fu_1714_p2);

assign xor_ln88_25_fu_2006_p2 = (and_ln88_22_fu_1994_p2 ^ and_ln87_22_fu_1940_p2);

assign xor_ln88_26_fu_2012_p2 = (and_ln88_23_fu_2000_p2 ^ and_ln88_20_fu_1982_p2);

assign xor_ln88_27_fu_2018_p2 = (xor_ln88_26_fu_2012_p2 ^ and_ln88_21_fu_1988_p2);

assign xor_ln88_28_fu_2024_p2 = (xor_ln88_27_fu_2018_p2 ^ xor_ln88_25_fu_2006_p2);

assign xor_ln88_29_fu_2030_p2 = (xor_ln88_28_fu_2024_p2 ^ xor_ln87_28_fu_1970_p2);

assign xor_ln88_2_fu_402_p2 = (and_ln88_3_fu_384_p2 ^ and_ln87_2_fu_324_p2);

assign xor_ln88_30_fu_2386_p2 = (and_ln88_26_fu_2374_p2 ^ and_ln88_25_fu_2368_p2);

assign xor_ln88_31_fu_2392_p2 = (xor_ln88_30_fu_2386_p2 ^ and_ln88_24_fu_2362_p2);

assign xor_ln88_32_fu_2398_p2 = (and_ln88_27_fu_2380_p2 ^ and_ln87_26_fu_2320_p2);

assign xor_ln88_33_fu_2404_p2 = (xor_ln88_32_fu_2398_p2 ^ xor_ln87_32_fu_2344_p2);

assign xor_ln88_34_fu_2410_p2 = (xor_ln88_33_fu_2404_p2 ^ xor_ln88_31_fu_2392_p2);

assign xor_ln88_35_fu_2688_p2 = (and_ln88_30_fu_2676_p2 ^ and_ln88_29_fu_2670_p2);

assign xor_ln88_36_fu_2694_p2 = (xor_ln88_35_fu_2688_p2 ^ and_ln88_28_fu_2664_p2);

assign xor_ln88_37_fu_2700_p2 = (and_ln88_31_fu_2682_p2 ^ and_ln87_30_fu_2622_p2);

assign xor_ln88_38_fu_2706_p2 = (xor_ln88_37_fu_2700_p2 ^ xor_ln87_37_fu_2646_p2);

assign xor_ln88_39_fu_2712_p2 = (xor_ln88_38_fu_2706_p2 ^ xor_ln88_36_fu_2694_p2);

assign xor_ln88_3_fu_408_p2 = (xor_ln88_2_fu_402_p2 ^ xor_ln87_2_fu_348_p2);

assign xor_ln88_40_fu_2986_p2 = (and_ln88_34_fu_2974_p2 ^ and_ln87_34_fu_2920_p2);

assign xor_ln88_41_fu_2992_p2 = (and_ln88_35_fu_2980_p2 ^ and_ln88_32_fu_2962_p2);

assign xor_ln88_42_fu_2998_p2 = (xor_ln88_41_fu_2992_p2 ^ and_ln88_33_fu_2968_p2);

assign xor_ln88_43_fu_3004_p2 = (xor_ln88_42_fu_2998_p2 ^ xor_ln88_40_fu_2986_p2);

assign xor_ln88_44_fu_3010_p2 = (xor_ln88_43_fu_3004_p2 ^ xor_ln87_43_fu_2950_p2);

assign xor_ln88_45_fu_3592_p2 = (and_ln88_38_fu_3580_p2 ^ and_ln88_37_fu_3574_p2);

assign xor_ln88_46_fu_3598_p2 = (xor_ln88_45_fu_3592_p2 ^ and_ln88_36_fu_3568_p2);

assign xor_ln88_47_fu_3604_p2 = (and_ln88_39_fu_3586_p2 ^ and_ln87_38_fu_3526_p2);

assign xor_ln88_48_fu_3610_p2 = (xor_ln88_47_fu_3604_p2 ^ xor_ln87_47_fu_3550_p2);

assign xor_ln88_49_fu_3616_p2 = (xor_ln88_48_fu_3610_p2 ^ xor_ln88_46_fu_3598_p2);

assign xor_ln88_4_fu_414_p2 = (xor_ln88_3_fu_408_p2 ^ xor_ln88_1_fu_396_p2);

assign xor_ln88_50_fu_3894_p2 = (and_ln88_42_fu_3882_p2 ^ and_ln88_41_fu_3876_p2);

assign xor_ln88_51_fu_3900_p2 = (xor_ln88_50_fu_3894_p2 ^ and_ln88_40_fu_3870_p2);

assign xor_ln88_52_fu_3906_p2 = (and_ln88_43_fu_3888_p2 ^ and_ln87_42_fu_3828_p2);

assign xor_ln88_53_fu_3912_p2 = (xor_ln88_52_fu_3906_p2 ^ xor_ln87_52_fu_3852_p2);

assign xor_ln88_54_fu_3918_p2 = (xor_ln88_53_fu_3912_p2 ^ xor_ln88_51_fu_3900_p2);

assign xor_ln88_55_fu_4192_p2 = (and_ln88_46_fu_4180_p2 ^ and_ln87_46_fu_4126_p2);

assign xor_ln88_56_fu_4198_p2 = (and_ln88_47_fu_4186_p2 ^ and_ln88_44_fu_4168_p2);

assign xor_ln88_57_fu_4204_p2 = (xor_ln88_56_fu_4198_p2 ^ and_ln88_45_fu_4174_p2);

assign xor_ln88_58_fu_4210_p2 = (xor_ln88_57_fu_4204_p2 ^ xor_ln88_55_fu_4192_p2);

assign xor_ln88_59_fu_4216_p2 = (xor_ln88_58_fu_4210_p2 ^ xor_ln87_58_fu_4156_p2);

assign xor_ln88_5_fu_692_p2 = (and_ln88_6_fu_680_p2 ^ and_ln88_5_fu_674_p2);

assign xor_ln88_60_fu_4596_p2 = (and_ln88_50_fu_4584_p2 ^ and_ln88_49_fu_4578_p2);

assign xor_ln88_61_fu_4602_p2 = (xor_ln88_60_fu_4596_p2 ^ and_ln88_48_fu_4572_p2);

assign xor_ln88_62_fu_4608_p2 = (and_ln88_51_fu_4590_p2 ^ and_ln87_50_fu_4530_p2);

assign xor_ln88_63_fu_4614_p2 = (xor_ln88_62_fu_4608_p2 ^ xor_ln87_62_fu_4554_p2);

assign xor_ln88_64_fu_4620_p2 = (xor_ln88_63_fu_4614_p2 ^ xor_ln88_61_fu_4602_p2);

assign xor_ln88_65_fu_4910_p2 = (and_ln88_54_fu_4898_p2 ^ and_ln88_53_fu_4892_p2);

assign xor_ln88_66_fu_4916_p2 = (xor_ln88_65_fu_4910_p2 ^ and_ln88_52_fu_4886_p2);

assign xor_ln88_67_fu_4922_p2 = (and_ln88_55_fu_4904_p2 ^ and_ln87_54_fu_4844_p2);

assign xor_ln88_68_fu_4928_p2 = (xor_ln88_67_fu_4922_p2 ^ xor_ln87_67_fu_4868_p2);

assign xor_ln88_69_fu_4934_p2 = (xor_ln88_68_fu_4928_p2 ^ xor_ln88_66_fu_4916_p2);

assign xor_ln88_6_fu_698_p2 = (xor_ln88_5_fu_692_p2 ^ and_ln88_4_fu_668_p2);

assign xor_ln88_70_fu_5208_p2 = (and_ln88_58_fu_5196_p2 ^ and_ln87_58_fu_5142_p2);

assign xor_ln88_71_fu_5214_p2 = (and_ln88_59_fu_5202_p2 ^ and_ln88_56_fu_5184_p2);

assign xor_ln88_72_fu_5220_p2 = (xor_ln88_71_fu_5214_p2 ^ and_ln88_57_fu_5190_p2);

assign xor_ln88_73_fu_5226_p2 = (xor_ln88_72_fu_5220_p2 ^ xor_ln88_70_fu_5208_p2);

assign xor_ln88_74_fu_5232_p2 = (xor_ln88_73_fu_5226_p2 ^ xor_ln87_73_fu_5172_p2);

assign xor_ln88_75_fu_5588_p2 = (and_ln88_62_fu_5576_p2 ^ and_ln88_61_fu_5570_p2);

assign xor_ln88_76_fu_5594_p2 = (xor_ln88_75_fu_5588_p2 ^ and_ln88_60_fu_5564_p2);

assign xor_ln88_77_fu_5600_p2 = (and_ln88_63_fu_5582_p2 ^ and_ln87_62_fu_5522_p2);

assign xor_ln88_78_fu_5606_p2 = (xor_ln88_77_fu_5600_p2 ^ xor_ln87_77_fu_5546_p2);

assign xor_ln88_79_fu_5612_p2 = (xor_ln88_78_fu_5606_p2 ^ xor_ln88_76_fu_5594_p2);

assign xor_ln88_7_fu_704_p2 = (and_ln88_7_fu_686_p2 ^ and_ln87_6_fu_626_p2);

assign xor_ln88_80_fu_5890_p2 = (and_ln88_66_fu_5878_p2 ^ and_ln88_65_fu_5872_p2);

assign xor_ln88_81_fu_5896_p2 = (xor_ln88_80_fu_5890_p2 ^ and_ln88_64_fu_5866_p2);

assign xor_ln88_82_fu_5902_p2 = (and_ln88_67_fu_5884_p2 ^ and_ln87_66_fu_5824_p2);

assign xor_ln88_83_fu_5908_p2 = (xor_ln88_82_fu_5902_p2 ^ xor_ln87_82_fu_5848_p2);

assign xor_ln88_84_fu_5914_p2 = (xor_ln88_83_fu_5908_p2 ^ xor_ln88_81_fu_5896_p2);

assign xor_ln88_85_fu_6188_p2 = (and_ln88_70_fu_6176_p2 ^ and_ln87_70_fu_6122_p2);

assign xor_ln88_86_fu_6194_p2 = (and_ln88_71_fu_6182_p2 ^ and_ln88_68_fu_6164_p2);

assign xor_ln88_87_fu_6200_p2 = (xor_ln88_86_fu_6194_p2 ^ and_ln88_69_fu_6170_p2);

assign xor_ln88_88_fu_6206_p2 = (xor_ln88_87_fu_6200_p2 ^ xor_ln88_85_fu_6188_p2);

assign xor_ln88_89_fu_6212_p2 = (xor_ln88_88_fu_6206_p2 ^ xor_ln87_88_fu_6152_p2);

assign xor_ln88_8_fu_710_p2 = (xor_ln88_7_fu_704_p2 ^ xor_ln87_7_fu_650_p2);

assign xor_ln88_90_fu_6726_p2 = (and_ln88_74_fu_6714_p2 ^ and_ln88_73_fu_6708_p2);

assign xor_ln88_91_fu_6732_p2 = (xor_ln88_90_fu_6726_p2 ^ and_ln88_72_fu_6702_p2);

assign xor_ln88_92_fu_6738_p2 = (and_ln88_75_fu_6720_p2 ^ and_ln87_74_fu_6660_p2);

assign xor_ln88_93_fu_6744_p2 = (xor_ln88_92_fu_6738_p2 ^ xor_ln87_92_fu_6684_p2);

assign xor_ln88_94_fu_6750_p2 = (xor_ln88_93_fu_6744_p2 ^ xor_ln88_91_fu_6732_p2);

assign xor_ln88_95_fu_7028_p2 = (and_ln88_78_fu_7016_p2 ^ and_ln88_77_fu_7010_p2);

assign xor_ln88_96_fu_7034_p2 = (xor_ln88_95_fu_7028_p2 ^ and_ln88_76_fu_7004_p2);

assign xor_ln88_97_fu_7040_p2 = (and_ln88_79_fu_7022_p2 ^ and_ln87_78_fu_6962_p2);

assign xor_ln88_98_fu_7046_p2 = (xor_ln88_97_fu_7040_p2 ^ xor_ln87_97_fu_6986_p2);

assign xor_ln88_99_fu_7052_p2 = (xor_ln88_98_fu_7046_p2 ^ xor_ln88_96_fu_7034_p2);

assign xor_ln88_9_fu_716_p2 = (xor_ln88_8_fu_710_p2 ^ xor_ln88_6_fu_698_p2);

assign xor_ln88_fu_390_p2 = (and_ln88_2_fu_378_p2 ^ and_ln88_1_fu_372_p2);

assign xor_ln91_100_fu_3966_p2 = (and_ln87_42_fu_3828_p2 ^ and_ln86_42_fu_3770_p2);

assign xor_ln91_101_fu_3972_p2 = (and_ln88_43_fu_3888_p2 ^ and_ln87_43_fu_3834_p2);

assign xor_ln91_102_fu_3978_p2 = (xor_ln91_101_fu_3972_p2 ^ and_ln91_10_fu_3942_p2);

assign xor_ln91_103_fu_3984_p2 = (xor_ln91_102_fu_3978_p2 ^ xor_ln91_100_fu_3966_p2);

assign xor_ln91_104_fu_4246_p2 = (and_ln91_11_fu_4240_p2 ^ and_ln88_47_fu_4186_p2);

assign xor_ln91_105_fu_4252_p2 = (and_ln87_46_fu_4126_p2 ^ and_ln86_46_fu_4068_p2);

assign xor_ln91_106_fu_4258_p2 = (xor_ln91_105_fu_4252_p2 ^ xor_ln91_104_fu_4246_p2);

assign xor_ln91_107_fu_4264_p2 = (and_ln90_34_fu_4228_p2 ^ and_ln90_33_fu_4222_p2);

assign xor_ln91_108_fu_4270_p2 = (and_ln88_45_fu_4174_p2 ^ and_ln87_47_fu_4150_p2);

assign xor_ln91_109_fu_4276_p2 = (xor_ln91_108_fu_4270_p2 ^ and_ln90_35_fu_4234_p2);

assign xor_ln91_10_fu_474_p2 = (xor_ln91_8_fu_468_p2 ^ and_ln91_fu_438_p2);

assign xor_ln91_110_fu_4282_p2 = (xor_ln91_109_fu_4276_p2 ^ xor_ln91_107_fu_4264_p2);

assign xor_ln91_111_fu_4650_p2 = (and_ln90_37_fu_4632_p2 ^ and_ln90_36_fu_4626_p2);

assign xor_ln91_112_fu_4656_p2 = (and_ln90_38_fu_4638_p2 ^ and_ln88_49_fu_4578_p2);

assign xor_ln91_113_fu_4662_p2 = (xor_ln91_112_fu_4656_p2 ^ xor_ln91_111_fu_4650_p2);

assign xor_ln91_114_fu_4668_p2 = (and_ln87_50_fu_4530_p2 ^ and_ln86_50_fu_4472_p2);

assign xor_ln91_115_fu_4674_p2 = (and_ln88_51_fu_4590_p2 ^ and_ln87_51_fu_4536_p2);

assign xor_ln91_116_fu_4680_p2 = (xor_ln91_115_fu_4674_p2 ^ and_ln91_12_fu_4644_p2);

assign xor_ln91_117_fu_4686_p2 = (xor_ln91_116_fu_4680_p2 ^ xor_ln91_114_fu_4668_p2);

assign xor_ln91_118_fu_4964_p2 = (and_ln90_40_fu_4946_p2 ^ and_ln90_39_fu_4940_p2);

assign xor_ln91_119_fu_4970_p2 = (and_ln90_41_fu_4952_p2 ^ and_ln88_53_fu_4892_p2);

assign xor_ln91_11_fu_2102_p2 = (xor_ln91_68_fu_2096_p2 ^ xor_ln91_64_fu_2072_p2);

assign xor_ln91_120_fu_4976_p2 = (xor_ln91_119_fu_4970_p2 ^ xor_ln91_118_fu_4964_p2);

assign xor_ln91_121_fu_4982_p2 = (and_ln87_54_fu_4844_p2 ^ and_ln86_54_fu_4786_p2);

assign xor_ln91_122_fu_4988_p2 = (and_ln88_55_fu_4904_p2 ^ and_ln87_55_fu_4850_p2);

assign xor_ln91_123_fu_4994_p2 = (xor_ln91_122_fu_4988_p2 ^ and_ln91_13_fu_4958_p2);

assign xor_ln91_124_fu_5000_p2 = (xor_ln91_123_fu_4994_p2 ^ xor_ln91_121_fu_4982_p2);

assign xor_ln91_125_fu_5262_p2 = (and_ln91_14_fu_5256_p2 ^ and_ln88_59_fu_5202_p2);

assign xor_ln91_126_fu_5268_p2 = (and_ln87_58_fu_5142_p2 ^ and_ln86_58_fu_5084_p2);

assign xor_ln91_127_fu_5274_p2 = (xor_ln91_126_fu_5268_p2 ^ xor_ln91_125_fu_5262_p2);

assign xor_ln91_128_fu_5280_p2 = (and_ln90_43_fu_5244_p2 ^ and_ln90_42_fu_5238_p2);

assign xor_ln91_129_fu_5286_p2 = (and_ln88_57_fu_5190_p2 ^ and_ln87_59_fu_5166_p2);

assign xor_ln91_12_fu_480_p2 = (xor_ln91_6_fu_462_p2 ^ xor_ln91_10_fu_474_p2);

assign xor_ln91_130_fu_5292_p2 = (xor_ln91_129_fu_5286_p2 ^ and_ln90_44_fu_5250_p2);

assign xor_ln91_131_fu_5298_p2 = (xor_ln91_130_fu_5292_p2 ^ xor_ln91_128_fu_5280_p2);

assign xor_ln91_132_fu_5642_p2 = (and_ln90_46_fu_5624_p2 ^ and_ln90_45_fu_5618_p2);

assign xor_ln91_133_fu_5648_p2 = (and_ln90_47_fu_5630_p2 ^ and_ln88_61_fu_5570_p2);

assign xor_ln91_134_fu_5654_p2 = (xor_ln91_133_fu_5648_p2 ^ xor_ln91_132_fu_5642_p2);

assign xor_ln91_135_fu_5660_p2 = (and_ln87_62_fu_5522_p2 ^ and_ln86_62_fu_5464_p2);

assign xor_ln91_136_fu_5666_p2 = (and_ln88_63_fu_5582_p2 ^ and_ln87_63_fu_5528_p2);

assign xor_ln91_137_fu_5672_p2 = (xor_ln91_136_fu_5666_p2 ^ and_ln91_15_fu_5636_p2);

assign xor_ln91_138_fu_5678_p2 = (xor_ln91_137_fu_5672_p2 ^ xor_ln91_135_fu_5660_p2);

assign xor_ln91_139_fu_5944_p2 = (and_ln90_49_fu_5926_p2 ^ and_ln90_48_fu_5920_p2);

assign xor_ln91_13_fu_2482_p2 = (xor_ln91_75_fu_2476_p2 ^ xor_ln91_71_fu_2452_p2);

assign xor_ln91_140_fu_5950_p2 = (and_ln90_50_fu_5932_p2 ^ and_ln88_65_fu_5872_p2);

assign xor_ln91_141_fu_5956_p2 = (xor_ln91_140_fu_5950_p2 ^ xor_ln91_139_fu_5944_p2);

assign xor_ln91_142_fu_5962_p2 = (and_ln87_66_fu_5824_p2 ^ and_ln86_66_fu_5766_p2);

assign xor_ln91_143_fu_5968_p2 = (and_ln88_67_fu_5884_p2 ^ and_ln87_67_fu_5830_p2);

assign xor_ln91_144_fu_5974_p2 = (xor_ln91_143_fu_5968_p2 ^ and_ln91_16_fu_5938_p2);

assign xor_ln91_145_fu_5980_p2 = (xor_ln91_144_fu_5974_p2 ^ xor_ln91_142_fu_5962_p2);

assign xor_ln91_146_fu_6242_p2 = (and_ln91_17_fu_6236_p2 ^ and_ln88_71_fu_6182_p2);

assign xor_ln91_147_fu_6248_p2 = (and_ln87_70_fu_6122_p2 ^ and_ln86_70_fu_6064_p2);

assign xor_ln91_148_fu_6254_p2 = (xor_ln91_147_fu_6248_p2 ^ xor_ln91_146_fu_6242_p2);

assign xor_ln91_149_fu_6260_p2 = (and_ln90_52_fu_6224_p2 ^ and_ln90_51_fu_6218_p2);

assign xor_ln91_14_fu_746_p2 = (and_ln90_4_fu_728_p2 ^ and_ln90_3_fu_722_p2);

assign xor_ln91_150_fu_6266_p2 = (and_ln88_69_fu_6170_p2 ^ and_ln87_71_fu_6146_p2);

assign xor_ln91_151_fu_6272_p2 = (xor_ln91_150_fu_6266_p2 ^ and_ln90_53_fu_6230_p2);

assign xor_ln91_152_fu_6278_p2 = (xor_ln91_151_fu_6272_p2 ^ xor_ln91_149_fu_6260_p2);

assign xor_ln91_153_fu_6780_p2 = (and_ln90_55_fu_6762_p2 ^ and_ln90_54_fu_6756_p2);

assign xor_ln91_154_fu_6786_p2 = (and_ln90_56_fu_6768_p2 ^ and_ln88_73_fu_6708_p2);

assign xor_ln91_155_fu_6792_p2 = (xor_ln91_154_fu_6786_p2 ^ xor_ln91_153_fu_6780_p2);

assign xor_ln91_156_fu_6798_p2 = (and_ln87_74_fu_6660_p2 ^ and_ln86_74_fu_6602_p2);

assign xor_ln91_157_fu_6804_p2 = (and_ln88_75_fu_6720_p2 ^ and_ln87_75_fu_6666_p2);

assign xor_ln91_158_fu_6810_p2 = (xor_ln91_157_fu_6804_p2 ^ and_ln91_18_fu_6774_p2);

assign xor_ln91_159_fu_6816_p2 = (xor_ln91_158_fu_6810_p2 ^ xor_ln91_156_fu_6798_p2);

assign xor_ln91_15_fu_2784_p2 = (xor_ln91_82_fu_2778_p2 ^ xor_ln91_78_fu_2754_p2);

assign xor_ln91_160_fu_7082_p2 = (and_ln90_58_fu_7064_p2 ^ and_ln90_57_fu_7058_p2);

assign xor_ln91_161_fu_7088_p2 = (and_ln90_59_fu_7070_p2 ^ and_ln88_77_fu_7010_p2);

assign xor_ln91_162_fu_7094_p2 = (xor_ln91_161_fu_7088_p2 ^ xor_ln91_160_fu_7082_p2);

assign xor_ln91_163_fu_7100_p2 = (and_ln87_78_fu_6962_p2 ^ and_ln86_78_fu_6904_p2);

assign xor_ln91_164_fu_7106_p2 = (and_ln88_79_fu_7022_p2 ^ and_ln87_79_fu_6968_p2);

assign xor_ln91_165_fu_7112_p2 = (xor_ln91_164_fu_7106_p2 ^ and_ln91_19_fu_7076_p2);

assign xor_ln91_166_fu_7118_p2 = (xor_ln91_165_fu_7112_p2 ^ xor_ln91_163_fu_7100_p2);

assign xor_ln91_167_fu_7380_p2 = (and_ln91_20_fu_7374_p2 ^ and_ln88_83_fu_7320_p2);

assign xor_ln91_168_fu_7386_p2 = (and_ln87_82_fu_7260_p2 ^ and_ln86_82_fu_7202_p2);

assign xor_ln91_169_fu_7392_p2 = (xor_ln91_168_fu_7386_p2 ^ xor_ln91_167_fu_7380_p2);

assign xor_ln91_16_fu_752_p2 = (and_ln90_5_fu_734_p2 ^ and_ln88_5_fu_674_p2);

assign xor_ln91_170_fu_7398_p2 = (and_ln90_61_fu_7362_p2 ^ and_ln90_60_fu_7356_p2);

assign xor_ln91_171_fu_7404_p2 = (and_ln88_81_fu_7308_p2 ^ and_ln87_83_fu_7284_p2);

assign xor_ln91_172_fu_7410_p2 = (xor_ln91_171_fu_7404_p2 ^ and_ln90_62_fu_7368_p2);

assign xor_ln91_173_fu_7416_p2 = (xor_ln91_172_fu_7410_p2 ^ xor_ln91_170_fu_7398_p2);

assign xor_ln91_174_fu_7784_p2 = (and_ln90_64_fu_7766_p2 ^ and_ln90_63_fu_7760_p2);

assign xor_ln91_175_fu_7790_p2 = (and_ln90_65_fu_7772_p2 ^ and_ln88_85_fu_7712_p2);

assign xor_ln91_176_fu_7796_p2 = (xor_ln91_175_fu_7790_p2 ^ xor_ln91_174_fu_7784_p2);

assign xor_ln91_177_fu_7802_p2 = (and_ln87_86_fu_7664_p2 ^ and_ln86_86_fu_7606_p2);

assign xor_ln91_178_fu_7808_p2 = (and_ln88_87_fu_7724_p2 ^ and_ln87_87_fu_7670_p2);

assign xor_ln91_179_fu_7814_p2 = (xor_ln91_178_fu_7808_p2 ^ and_ln91_21_fu_7778_p2);

assign xor_ln91_17_fu_3082_p2 = (xor_ln91_89_fu_3076_p2 ^ xor_ln91_85_fu_3052_p2);

assign xor_ln91_180_fu_7820_p2 = (xor_ln91_179_fu_7814_p2 ^ xor_ln91_177_fu_7802_p2);

assign xor_ln91_181_fu_8098_p2 = (and_ln90_67_fu_8080_p2 ^ and_ln90_66_fu_8074_p2);

assign xor_ln91_182_fu_8104_p2 = (and_ln90_68_fu_8086_p2 ^ and_ln88_89_fu_8026_p2);

assign xor_ln91_183_fu_8110_p2 = (xor_ln91_182_fu_8104_p2 ^ xor_ln91_181_fu_8098_p2);

assign xor_ln91_184_fu_8116_p2 = (and_ln87_90_fu_7978_p2 ^ and_ln86_90_fu_7920_p2);

assign xor_ln91_185_fu_8122_p2 = (and_ln88_91_fu_8038_p2 ^ and_ln87_91_fu_7984_p2);

assign xor_ln91_186_fu_8128_p2 = (xor_ln91_185_fu_8122_p2 ^ and_ln91_22_fu_8092_p2);

assign xor_ln91_187_fu_8134_p2 = (xor_ln91_186_fu_8128_p2 ^ xor_ln91_184_fu_8116_p2);

assign xor_ln91_188_fu_8396_p2 = (and_ln91_23_fu_8390_p2 ^ and_ln88_95_fu_8336_p2);

assign xor_ln91_189_fu_8402_p2 = (and_ln87_94_fu_8276_p2 ^ and_ln86_94_fu_8218_p2);

assign xor_ln91_18_fu_758_p2 = (xor_ln91_16_fu_752_p2 ^ xor_ln91_14_fu_746_p2);

assign xor_ln91_190_fu_8408_p2 = (xor_ln91_189_fu_8402_p2 ^ xor_ln91_188_fu_8396_p2);

assign xor_ln91_191_fu_8414_p2 = (and_ln90_70_fu_8378_p2 ^ and_ln90_69_fu_8372_p2);

assign xor_ln91_192_fu_8420_p2 = (and_ln88_93_fu_8324_p2 ^ and_ln87_95_fu_8300_p2);

assign xor_ln91_193_fu_8426_p2 = (xor_ln91_192_fu_8420_p2 ^ and_ln90_71_fu_8384_p2);

assign xor_ln91_194_fu_8432_p2 = (xor_ln91_193_fu_8426_p2 ^ xor_ln91_191_fu_8414_p2);

assign xor_ln91_195_fu_8776_p2 = (and_ln90_73_fu_8758_p2 ^ and_ln90_72_fu_8752_p2);

assign xor_ln91_196_fu_8782_p2 = (and_ln90_74_fu_8764_p2 ^ and_ln88_97_fu_8704_p2);

assign xor_ln91_197_fu_8788_p2 = (xor_ln91_196_fu_8782_p2 ^ xor_ln91_195_fu_8776_p2);

assign xor_ln91_198_fu_8794_p2 = (and_ln87_98_fu_8656_p2 ^ and_ln86_98_fu_8598_p2);

assign xor_ln91_199_fu_8800_p2 = (and_ln88_99_fu_8716_p2 ^ and_ln87_99_fu_8662_p2);

assign xor_ln91_19_fu_3688_p2 = (xor_ln91_96_fu_3682_p2 ^ xor_ln91_92_fu_3658_p2);

assign xor_ln91_1_fu_486_p2 = (xor_ln91_4_fu_456_p2 ^ xor_ln91_12_fu_480_p2);

assign xor_ln91_200_fu_8806_p2 = (xor_ln91_199_fu_8800_p2 ^ and_ln91_24_fu_8770_p2);

assign xor_ln91_201_fu_8812_p2 = (xor_ln91_200_fu_8806_p2 ^ xor_ln91_198_fu_8794_p2);

assign xor_ln91_202_fu_9078_p2 = (and_ln90_76_fu_9060_p2 ^ and_ln90_75_fu_9054_p2);

assign xor_ln91_203_fu_9084_p2 = (and_ln90_77_fu_9066_p2 ^ and_ln88_101_fu_9006_p2);

assign xor_ln91_204_fu_9090_p2 = (xor_ln91_203_fu_9084_p2 ^ xor_ln91_202_fu_9078_p2);

assign xor_ln91_205_fu_9096_p2 = (and_ln87_102_fu_8958_p2 ^ and_ln86_102_fu_8900_p2);

assign xor_ln91_206_fu_9102_p2 = (and_ln88_103_fu_9018_p2 ^ and_ln87_103_fu_8964_p2);

assign xor_ln91_207_fu_9108_p2 = (xor_ln91_206_fu_9102_p2 ^ and_ln91_25_fu_9072_p2);

assign xor_ln91_208_fu_9114_p2 = (xor_ln91_207_fu_9108_p2 ^ xor_ln91_205_fu_9096_p2);

assign xor_ln91_209_fu_9376_p2 = (and_ln91_26_fu_9370_p2 ^ and_ln88_107_fu_9316_p2);

assign xor_ln91_20_fu_764_p2 = (and_ln87_6_fu_626_p2 ^ and_ln86_6_fu_568_p2);

assign xor_ln91_210_fu_9382_p2 = (and_ln87_106_fu_9256_p2 ^ and_ln86_106_fu_9198_p2);

assign xor_ln91_211_fu_9388_p2 = (xor_ln91_210_fu_9382_p2 ^ xor_ln91_209_fu_9376_p2);

assign xor_ln91_212_fu_9394_p2 = (and_ln90_79_fu_9358_p2 ^ and_ln90_78_fu_9352_p2);

assign xor_ln91_213_fu_9400_p2 = (and_ln88_105_fu_9304_p2 ^ and_ln87_107_fu_9280_p2);

assign xor_ln91_214_fu_9406_p2 = (xor_ln91_213_fu_9400_p2 ^ and_ln90_80_fu_9364_p2);

assign xor_ln91_215_fu_9412_p2 = (xor_ln91_214_fu_9406_p2 ^ xor_ln91_212_fu_9394_p2);

assign xor_ln91_21_fu_3990_p2 = (xor_ln91_99_fu_3960_p2 ^ xor_ln91_103_fu_3984_p2);

assign xor_ln91_22_fu_770_p2 = (and_ln88_7_fu_686_p2 ^ and_ln87_7_fu_632_p2);

assign xor_ln91_23_fu_4288_p2 = (xor_ln91_110_fu_4282_p2 ^ xor_ln91_106_fu_4258_p2);

assign xor_ln91_24_fu_776_p2 = (xor_ln91_22_fu_770_p2 ^ and_ln91_1_fu_740_p2);

assign xor_ln91_25_fu_4692_p2 = (xor_ln91_117_fu_4686_p2 ^ xor_ln91_113_fu_4662_p2);

assign xor_ln91_26_fu_782_p2 = (xor_ln91_24_fu_776_p2 ^ xor_ln91_20_fu_764_p2);

assign xor_ln91_27_fu_5006_p2 = (xor_ln91_124_fu_5000_p2 ^ xor_ln91_120_fu_4976_p2);

assign xor_ln91_28_fu_1044_p2 = (and_ln91_2_fu_1038_p2 ^ and_ln88_11_fu_984_p2);

assign xor_ln91_29_fu_5304_p2 = (xor_ln91_131_fu_5298_p2 ^ xor_ln91_127_fu_5274_p2);

assign xor_ln91_2_fu_450_p2 = (and_ln90_2_fu_432_p2 ^ and_ln88_1_fu_372_p2);

assign xor_ln91_30_fu_1050_p2 = (and_ln87_10_fu_924_p2 ^ and_ln86_10_fu_866_p2);

assign xor_ln91_31_fu_5684_p2 = (xor_ln91_138_fu_5678_p2 ^ xor_ln91_134_fu_5654_p2);

assign xor_ln91_32_fu_1056_p2 = (xor_ln91_30_fu_1050_p2 ^ xor_ln91_28_fu_1044_p2);

assign xor_ln91_33_fu_5986_p2 = (xor_ln91_145_fu_5980_p2 ^ xor_ln91_141_fu_5956_p2);

assign xor_ln91_34_fu_1062_p2 = (and_ln90_7_fu_1026_p2 ^ and_ln90_6_fu_1020_p2);

assign xor_ln91_35_fu_6284_p2 = (xor_ln91_152_fu_6278_p2 ^ xor_ln91_148_fu_6254_p2);

assign xor_ln91_36_fu_1068_p2 = (and_ln88_9_fu_972_p2 ^ and_ln87_11_fu_948_p2);

assign xor_ln91_37_fu_6822_p2 = (xor_ln91_159_fu_6816_p2 ^ xor_ln91_155_fu_6792_p2);

assign xor_ln91_38_fu_1074_p2 = (xor_ln91_36_fu_1068_p2 ^ and_ln90_8_fu_1032_p2);

assign xor_ln91_39_fu_7124_p2 = (xor_ln91_166_fu_7118_p2 ^ xor_ln91_162_fu_7094_p2);

assign xor_ln91_3_fu_788_p2 = (xor_ln91_26_fu_782_p2 ^ xor_ln91_18_fu_758_p2);

assign xor_ln91_40_fu_1080_p2 = (xor_ln91_38_fu_1074_p2 ^ xor_ln91_34_fu_1062_p2);

assign xor_ln91_41_fu_7422_p2 = (xor_ln91_173_fu_7416_p2 ^ xor_ln91_169_fu_7392_p2);

assign xor_ln91_42_fu_1448_p2 = (and_ln90_9_fu_1424_p2 ^ and_ln90_10_fu_1430_p2);

assign xor_ln91_43_fu_7826_p2 = (xor_ln91_180_fu_7820_p2 ^ xor_ln91_176_fu_7796_p2);

assign xor_ln91_44_fu_1454_p2 = (and_ln90_11_fu_1436_p2 ^ and_ln88_13_fu_1376_p2);

assign xor_ln91_45_fu_8140_p2 = (xor_ln91_187_fu_8134_p2 ^ xor_ln91_183_fu_8110_p2);

assign xor_ln91_46_fu_1460_p2 = (xor_ln91_44_fu_1454_p2 ^ xor_ln91_42_fu_1448_p2);

assign xor_ln91_47_fu_8438_p2 = (xor_ln91_194_fu_8432_p2 ^ xor_ln91_190_fu_8408_p2);

assign xor_ln91_48_fu_1466_p2 = (and_ln87_14_fu_1328_p2 ^ and_ln86_14_fu_1270_p2);

assign xor_ln91_49_fu_8818_p2 = (xor_ln91_201_fu_8812_p2 ^ xor_ln91_197_fu_8788_p2);

assign xor_ln91_4_fu_456_p2 = (xor_ln91_fu_444_p2 ^ xor_ln91_2_fu_450_p2);

assign xor_ln91_50_fu_1472_p2 = (and_ln88_15_fu_1388_p2 ^ and_ln87_15_fu_1334_p2);

assign xor_ln91_51_fu_9120_p2 = (xor_ln91_208_fu_9114_p2 ^ xor_ln91_204_fu_9090_p2);

assign xor_ln91_52_fu_1478_p2 = (xor_ln91_50_fu_1472_p2 ^ and_ln91_3_fu_1442_p2);

assign xor_ln91_53_fu_9418_p2 = (xor_ln91_215_fu_9412_p2 ^ xor_ln91_211_fu_9388_p2);

assign xor_ln91_54_fu_1484_p2 = (xor_ln91_52_fu_1478_p2 ^ xor_ln91_48_fu_1466_p2);

assign xor_ln91_55_fu_1762_p2 = (and_ln90_13_fu_1744_p2 ^ and_ln90_12_fu_1738_p2);

assign xor_ln91_56_fu_1768_p2 = (and_ln90_14_fu_1750_p2 ^ and_ln88_17_fu_1690_p2);

assign xor_ln91_57_fu_1774_p2 = (xor_ln91_56_fu_1768_p2 ^ xor_ln91_55_fu_1762_p2);

assign xor_ln91_58_fu_1780_p2 = (and_ln87_18_fu_1642_p2 ^ and_ln86_18_fu_1584_p2);

assign xor_ln91_59_fu_1786_p2 = (and_ln88_19_fu_1702_p2 ^ and_ln87_19_fu_1648_p2);

assign xor_ln91_5_fu_1086_p2 = (xor_ln91_40_fu_1080_p2 ^ xor_ln91_32_fu_1056_p2);

assign xor_ln91_60_fu_1792_p2 = (xor_ln91_59_fu_1786_p2 ^ and_ln91_4_fu_1756_p2);

assign xor_ln91_61_fu_1798_p2 = (xor_ln91_60_fu_1792_p2 ^ xor_ln91_58_fu_1780_p2);

assign xor_ln91_62_fu_2060_p2 = (and_ln91_5_fu_2054_p2 ^ and_ln88_23_fu_2000_p2);

assign xor_ln91_63_fu_2066_p2 = (and_ln87_22_fu_1940_p2 ^ and_ln86_22_fu_1882_p2);

assign xor_ln91_64_fu_2072_p2 = (xor_ln91_63_fu_2066_p2 ^ xor_ln91_62_fu_2060_p2);

assign xor_ln91_65_fu_2078_p2 = (and_ln90_16_fu_2042_p2 ^ and_ln90_15_fu_2036_p2);

assign xor_ln91_66_fu_2084_p2 = (and_ln88_21_fu_1988_p2 ^ and_ln87_23_fu_1964_p2);

assign xor_ln91_67_fu_2090_p2 = (xor_ln91_66_fu_2084_p2 ^ and_ln90_17_fu_2048_p2);

assign xor_ln91_68_fu_2096_p2 = (xor_ln91_67_fu_2090_p2 ^ xor_ln91_65_fu_2078_p2);

assign xor_ln91_69_fu_2440_p2 = (and_ln90_19_fu_2422_p2 ^ and_ln90_18_fu_2416_p2);

assign xor_ln91_6_fu_462_p2 = (and_ln87_2_fu_324_p2 ^ and_ln86_2_fu_266_p2);

assign xor_ln91_70_fu_2446_p2 = (and_ln90_20_fu_2428_p2 ^ and_ln88_25_fu_2368_p2);

assign xor_ln91_71_fu_2452_p2 = (xor_ln91_70_fu_2446_p2 ^ xor_ln91_69_fu_2440_p2);

assign xor_ln91_72_fu_2458_p2 = (and_ln87_26_fu_2320_p2 ^ and_ln86_26_fu_2262_p2);

assign xor_ln91_73_fu_2464_p2 = (and_ln88_27_fu_2380_p2 ^ and_ln87_27_fu_2326_p2);

assign xor_ln91_74_fu_2470_p2 = (xor_ln91_73_fu_2464_p2 ^ and_ln91_6_fu_2434_p2);

assign xor_ln91_75_fu_2476_p2 = (xor_ln91_74_fu_2470_p2 ^ xor_ln91_72_fu_2458_p2);

assign xor_ln91_76_fu_2742_p2 = (and_ln90_22_fu_2724_p2 ^ and_ln90_21_fu_2718_p2);

assign xor_ln91_77_fu_2748_p2 = (and_ln90_23_fu_2730_p2 ^ and_ln88_29_fu_2670_p2);

assign xor_ln91_78_fu_2754_p2 = (xor_ln91_77_fu_2748_p2 ^ xor_ln91_76_fu_2742_p2);

assign xor_ln91_79_fu_2760_p2 = (and_ln87_30_fu_2622_p2 ^ and_ln86_30_fu_2564_p2);

assign xor_ln91_7_fu_1490_p2 = (xor_ln91_54_fu_1484_p2 ^ xor_ln91_46_fu_1460_p2);

assign xor_ln91_80_fu_2766_p2 = (and_ln88_31_fu_2682_p2 ^ and_ln87_31_fu_2628_p2);

assign xor_ln91_81_fu_2772_p2 = (xor_ln91_80_fu_2766_p2 ^ and_ln91_7_fu_2736_p2);

assign xor_ln91_82_fu_2778_p2 = (xor_ln91_81_fu_2772_p2 ^ xor_ln91_79_fu_2760_p2);

assign xor_ln91_83_fu_3040_p2 = (and_ln91_8_fu_3034_p2 ^ and_ln88_35_fu_2980_p2);

assign xor_ln91_84_fu_3046_p2 = (and_ln87_34_fu_2920_p2 ^ and_ln86_34_fu_2862_p2);

assign xor_ln91_85_fu_3052_p2 = (xor_ln91_84_fu_3046_p2 ^ xor_ln91_83_fu_3040_p2);

assign xor_ln91_86_fu_3058_p2 = (and_ln90_25_fu_3022_p2 ^ and_ln90_24_fu_3016_p2);

assign xor_ln91_87_fu_3064_p2 = (and_ln88_33_fu_2968_p2 ^ and_ln87_35_fu_2944_p2);

assign xor_ln91_88_fu_3070_p2 = (xor_ln91_87_fu_3064_p2 ^ and_ln90_26_fu_3028_p2);

assign xor_ln91_89_fu_3076_p2 = (xor_ln91_88_fu_3070_p2 ^ xor_ln91_86_fu_3058_p2);

assign xor_ln91_8_fu_468_p2 = (and_ln88_3_fu_384_p2 ^ and_ln87_3_fu_330_p2);

assign xor_ln91_90_fu_3646_p2 = (and_ln90_28_fu_3628_p2 ^ and_ln90_27_fu_3622_p2);

assign xor_ln91_91_fu_3652_p2 = (and_ln90_29_fu_3634_p2 ^ and_ln88_37_fu_3574_p2);

assign xor_ln91_92_fu_3658_p2 = (xor_ln91_91_fu_3652_p2 ^ xor_ln91_90_fu_3646_p2);

assign xor_ln91_93_fu_3664_p2 = (and_ln87_38_fu_3526_p2 ^ and_ln86_38_fu_3468_p2);

assign xor_ln91_94_fu_3670_p2 = (and_ln88_39_fu_3586_p2 ^ and_ln87_39_fu_3532_p2);

assign xor_ln91_95_fu_3676_p2 = (xor_ln91_94_fu_3670_p2 ^ and_ln91_9_fu_3640_p2);

assign xor_ln91_96_fu_3682_p2 = (xor_ln91_95_fu_3676_p2 ^ xor_ln91_93_fu_3664_p2);

assign xor_ln91_97_fu_3948_p2 = (and_ln90_31_fu_3930_p2 ^ and_ln90_30_fu_3924_p2);

assign xor_ln91_98_fu_3954_p2 = (and_ln90_32_fu_3936_p2 ^ and_ln88_41_fu_3876_p2);

assign xor_ln91_99_fu_3960_p2 = (xor_ln91_98_fu_3954_p2 ^ xor_ln91_97_fu_3948_p2);

assign xor_ln91_9_fu_1804_p2 = (xor_ln91_61_fu_1798_p2 ^ xor_ln91_57_fu_1774_p2);

assign xor_ln91_fu_444_p2 = (and_ln90_fu_420_p2 ^ and_ln90_1_fu_426_p2);

assign xor_ln99_14_fu_4710_p2 = (a1_17_fu_4400_p4 ^ a0_16_fu_3384_p2);

assign xor_ln99_16_fu_4722_p2 = (b1_17_fu_4410_p4 ^ b0_5_fu_3400_p2);

assign xor_ln99_24_fu_7844_p2 = (a1_21_fu_7534_p4 ^ a0_20_fu_7502_p4);

assign xor_ln99_26_fu_7856_p2 = (b1_21_fu_7544_p4 ^ b0_9_fu_7518_p4);

assign xor_ln99_4_fu_1520_p2 = (b1_13_fu_1208_p4 ^ b0_2_fu_200_p1);

assign xor_ln99_fu_1508_p2 = (a1_13_fu_1198_p4 ^ a0_13_fu_186_p1);

assign z0_10_fu_7494_p3 = {{xor_ln101_32_fu_7482_p2}, {xor_ln101_33_fu_7488_p2}};

assign z0_1_fu_1158_p3 = {{xor_ln101_2_fu_1146_p2}, {xor_ln101_3_fu_1152_p2}};

assign z0_4_fu_3292_p3 = {{xor_ln101_13_fu_3280_p2}, {xor_ln101_14_fu_3286_p2}};

assign z0_6_fu_4360_p3 = {{xor_ln101_17_fu_4348_p2}, {xor_ln101_18_fu_4354_p2}};

assign z1_11_fu_8510_p3 = {{xor_ln101_36_fu_8498_p2}, {xor_ln101_37_fu_8504_p2}};

assign z1_2_fu_2174_p3 = {{xor_ln101_6_fu_2162_p2}, {xor_ln101_7_fu_2168_p2}};

assign z1_6_fu_5376_p3 = {{xor_ln101_21_fu_5364_p2}, {xor_ln101_22_fu_5370_p2}};

assign z1_8_fu_6494_p3 = {{xor_ln101_28_fu_6482_p2}, {xor_ln101_29_fu_6488_p2}};

assign z2_4_fu_6350_p3 = {{xor_ln101_25_fu_6344_p2}, {xor_ln101_23_fu_6332_p2}};

assign z2_5_fu_9484_p3 = {{xor_ln101_40_fu_9478_p2}, {xor_ln101_38_fu_9466_p2}};

assign z2_6_fu_9622_p3 = {{a1_23_fu_9616_p2}, {a0_fu_9604_p2}};

assign z2_fu_3148_p3 = {{xor_ln101_10_fu_3142_p2}, {xor_ln101_8_fu_3130_p2}};

assign ap_return = {{xor_ln101_46_fu_9782_p2}, {xor_ln101_47_fu_9788_p2}};

endmodule //binary_tower_32b_mul
