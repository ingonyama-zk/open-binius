module binary_tower_32b_inv (
        ap_clk,
        ap_ce,
        ap_rst,
        a,
        ap_return
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;


input   ap_clk;
input   ap_ce;
input   ap_rst;
input  [31:0] a;
output  [31:0] ap_return;

wire   [0:0] a0_288_fu_244_p3;
reg   [0:0] a0_288_reg_13599;
(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] a0_288_reg_13599_pp0_iter1_reg;
wire   [0:0] a1_261_fu_252_p3;
reg   [0:0] a1_261_reg_13605;
reg   [0:0] a1_261_reg_13605_pp0_iter1_reg;
wire   [0:0] a0_339_fu_260_p2;
reg   [0:0] a0_339_reg_13610;
reg   [0:0] a0_339_reg_13610_pp0_iter1_reg;
wire   [0:0] a0_335_fu_362_p3;
reg   [0:0] a0_335_reg_13615;
reg   [0:0] a0_335_reg_13615_pp0_iter1_reg;
wire   [0:0] b0_3_fu_566_p2;
reg   [0:0] b0_3_reg_13623;
reg   [0:0] b0_3_reg_13623_pp0_iter1_reg;
wire   [0:0] b1_99_fu_572_p3;
reg   [0:0] b1_99_reg_13628;
reg   [0:0] b1_99_reg_13628_pp0_iter1_reg;
wire   [0:0] b_5_fu_592_p2;
reg   [0:0] b_5_reg_13633;
reg   [0:0] b_5_reg_13633_pp0_iter1_reg;
wire   [0:0] b0_5_fu_644_p3;
reg   [0:0] b0_5_reg_13638;
reg   [0:0] b0_5_reg_13638_pp0_iter1_reg;
wire   [0:0] b0_4_fu_672_p2;
reg   [0:0] b0_4_reg_13643;
reg   [0:0] b0_4_reg_13643_pp0_iter1_reg;
wire   [0:0] b1_100_fu_678_p3;
reg   [0:0] b1_100_reg_13648;
reg   [0:0] b1_100_reg_13648_pp0_iter1_reg;
wire   [0:0] b_9_fu_698_p2;
reg   [0:0] b_9_reg_13653;
reg   [0:0] b_9_reg_13653_pp0_iter1_reg;
wire   [0:0] b1_101_fu_744_p3;
reg   [0:0] b1_101_reg_13658;
reg   [0:0] b1_101_reg_13658_pp0_iter1_reg;
wire   [0:0] b_13_fu_764_p2;
reg   [0:0] b_13_reg_13663;
reg   [0:0] b_13_reg_13663_pp0_iter1_reg;
wire   [0:0] b0_11_fu_872_p3;
reg   [0:0] b0_11_reg_13668;
reg   [0:0] b0_11_reg_13668_pp0_iter1_reg;
wire   [0:0] b0_7_fu_942_p2;
reg   [0:0] b0_7_reg_13673;
reg   [0:0] b0_7_reg_13673_pp0_iter1_reg;
wire   [0:0] b1_103_fu_948_p3;
reg   [0:0] b1_103_reg_13678;
reg   [0:0] b1_103_reg_13678_pp0_iter1_reg;
wire   [0:0] b_18_fu_968_p2;
reg   [0:0] b_18_reg_13683;
reg   [0:0] b_18_reg_13683_pp0_iter1_reg;
wire   [0:0] b0_9_fu_1020_p3;
reg   [0:0] b0_9_reg_13688;
reg   [0:0] b0_9_reg_13688_pp0_iter1_reg;
wire   [0:0] b0_8_fu_1048_p2;
reg   [0:0] b0_8_reg_13693;
reg   [0:0] b0_8_reg_13693_pp0_iter1_reg;
wire   [0:0] b1_104_fu_1054_p3;
reg   [0:0] b1_104_reg_13698;
reg   [0:0] b1_104_reg_13698_pp0_iter1_reg;
wire   [0:0] b_22_fu_1074_p2;
reg   [0:0] b_22_reg_13703;
reg   [0:0] b_22_reg_13703_pp0_iter1_reg;
wire   [0:0] b1_105_fu_1120_p3;
reg   [0:0] b1_105_reg_13708;
reg   [0:0] b1_105_reg_13708_pp0_iter1_reg;
wire   [0:0] b_26_fu_1140_p2;
reg   [0:0] b_26_reg_13713;
reg   [0:0] b_26_reg_13713_pp0_iter1_reg;
wire   [0:0] b1_107_fu_1252_p3;
reg   [0:0] b1_107_reg_13718;
reg   [0:0] b1_107_reg_13718_pp0_iter1_reg;
wire   [0:0] b_31_fu_1272_p2;
reg   [0:0] b_31_reg_13723;
reg   [0:0] b_31_reg_13723_pp0_iter1_reg;
wire   [0:0] b0_13_fu_1324_p3;
reg   [0:0] b0_13_reg_13728;
reg   [0:0] b0_13_reg_13728_pp0_iter1_reg;
wire   [0:0] b0_12_fu_1352_p2;
reg   [0:0] b0_12_reg_13733;
reg   [0:0] b0_12_reg_13733_pp0_iter1_reg;
wire   [0:0] b1_108_fu_1358_p3;
reg   [0:0] b1_108_reg_13738;
reg   [0:0] b1_108_reg_13738_pp0_iter1_reg;
wire   [0:0] b_35_fu_1378_p2;
reg   [0:0] b_35_reg_13743;
reg   [0:0] b_35_reg_13743_pp0_iter1_reg;
wire   [0:0] b1_109_fu_1424_p3;
reg   [0:0] b1_109_reg_13748;
reg   [0:0] b1_109_reg_13748_pp0_iter1_reg;
wire   [0:0] b_39_fu_1444_p2;
reg   [0:0] b_39_reg_13753;
reg   [0:0] b_39_reg_13753_pp0_iter1_reg;
wire   [0:0] b0_29_fu_1674_p3;
reg   [0:0] b0_29_reg_13758;
reg   [0:0] b0_29_reg_13758_pp0_iter1_reg;
wire   [0:0] b0_16_fu_1802_p2;
reg   [0:0] b0_16_reg_13763;
reg   [0:0] b0_16_reg_13763_pp0_iter1_reg;
wire   [0:0] b1_112_fu_1808_p3;
reg   [0:0] b1_112_reg_13768;
reg   [0:0] b1_112_reg_13768_pp0_iter1_reg;
wire   [0:0] b_45_fu_1828_p2;
reg   [0:0] b_45_reg_13773;
reg   [0:0] b_45_reg_13773_pp0_iter1_reg;
wire   [0:0] b0_18_fu_1880_p3;
reg   [0:0] b0_18_reg_13778;
reg   [0:0] b0_18_reg_13778_pp0_iter1_reg;
wire   [0:0] b0_17_fu_1908_p2;
reg   [0:0] b0_17_reg_13783;
reg   [0:0] b0_17_reg_13783_pp0_iter1_reg;
wire   [0:0] b1_113_fu_1914_p3;
reg   [0:0] b1_113_reg_13788;
reg   [0:0] b1_113_reg_13788_pp0_iter1_reg;
wire   [0:0] b_49_fu_1934_p2;
reg   [0:0] b_49_reg_13793;
reg   [0:0] b_49_reg_13793_pp0_iter1_reg;
wire   [0:0] b1_114_fu_1980_p3;
reg   [0:0] b1_114_reg_13798;
reg   [0:0] b1_114_reg_13798_pp0_iter1_reg;
wire   [0:0] b_53_fu_2000_p2;
reg   [0:0] b_53_reg_13803;
reg   [0:0] b_53_reg_13803_pp0_iter1_reg;
wire   [0:0] b0_24_fu_2108_p3;
reg   [0:0] b0_24_reg_13808;
reg   [0:0] b0_24_reg_13808_pp0_iter1_reg;
wire   [0:0] b0_20_fu_2178_p2;
reg   [0:0] b0_20_reg_13813;
reg   [0:0] b0_20_reg_13813_pp0_iter1_reg;
wire   [0:0] b1_116_fu_2184_p3;
reg   [0:0] b1_116_reg_13818;
reg   [0:0] b1_116_reg_13818_pp0_iter1_reg;
wire   [0:0] b_58_fu_2204_p2;
reg   [0:0] b_58_reg_13823;
reg   [0:0] b_58_reg_13823_pp0_iter1_reg;
wire   [0:0] b0_22_fu_2256_p3;
reg   [0:0] b0_22_reg_13828;
reg   [0:0] b0_22_reg_13828_pp0_iter1_reg;
wire   [0:0] b0_21_fu_2284_p2;
reg   [0:0] b0_21_reg_13833;
reg   [0:0] b0_21_reg_13833_pp0_iter1_reg;
wire   [0:0] b1_117_fu_2290_p3;
reg   [0:0] b1_117_reg_13838;
reg   [0:0] b1_117_reg_13838_pp0_iter1_reg;
wire   [0:0] b_62_fu_2310_p2;
reg   [0:0] b_62_reg_13843;
reg   [0:0] b_62_reg_13843_pp0_iter1_reg;
wire   [0:0] b1_118_fu_2356_p3;
reg   [0:0] b1_118_reg_13848;
reg   [0:0] b1_118_reg_13848_pp0_iter1_reg;
wire   [0:0] b_66_fu_2376_p2;
reg   [0:0] b_66_reg_13853;
reg   [0:0] b_66_reg_13853_pp0_iter1_reg;
wire   [0:0] b1_120_fu_2488_p3;
reg   [0:0] b1_120_reg_13858;
reg   [0:0] b1_120_reg_13858_pp0_iter1_reg;
wire   [0:0] b_71_fu_2508_p2;
reg   [0:0] b_71_reg_13863;
reg   [0:0] b_71_reg_13863_pp0_iter1_reg;
wire   [0:0] b0_26_fu_2560_p3;
reg   [0:0] b0_26_reg_13868;
reg   [0:0] b0_26_reg_13868_pp0_iter1_reg;
wire   [0:0] b0_25_fu_2588_p2;
reg   [0:0] b0_25_reg_13873;
reg   [0:0] b0_25_reg_13873_pp0_iter1_reg;
wire   [0:0] b1_121_fu_2594_p3;
reg   [0:0] b1_121_reg_13878;
reg   [0:0] b1_121_reg_13878_pp0_iter1_reg;
wire   [0:0] b_75_fu_2614_p2;
reg   [0:0] b_75_reg_13883;
reg   [0:0] b_75_reg_13883_pp0_iter1_reg;
wire   [0:0] b1_122_fu_2660_p3;
reg   [0:0] b1_122_reg_13888;
reg   [0:0] b1_122_reg_13888_pp0_iter1_reg;
wire   [0:0] b_79_fu_2680_p2;
reg   [0:0] b_79_reg_13893;
reg   [0:0] b_79_reg_13893_pp0_iter1_reg;
wire   [0:0] b1_125_fu_2908_p3;
reg   [0:0] b1_125_reg_13898;
reg   [0:0] b1_125_reg_13898_pp0_iter1_reg;
wire   [0:0] b_85_fu_2928_p2;
reg   [0:0] b_85_reg_13903;
reg   [0:0] b_85_reg_13903_pp0_iter1_reg;
wire   [0:0] b0_31_fu_2980_p3;
reg   [0:0] b0_31_reg_13908;
reg   [0:0] b0_31_reg_13908_pp0_iter1_reg;
wire   [0:0] b0_30_fu_3008_p2;
reg   [0:0] b0_30_reg_13913;
reg   [0:0] b0_30_reg_13913_pp0_iter1_reg;
wire   [0:0] b1_126_fu_3014_p3;
reg   [0:0] b1_126_reg_13918;
reg   [0:0] b1_126_reg_13918_pp0_iter1_reg;
wire   [0:0] b_89_fu_3034_p2;
reg   [0:0] b_89_reg_13923;
reg   [0:0] b_89_reg_13923_pp0_iter1_reg;
wire   [0:0] b1_127_fu_3080_p3;
reg   [0:0] b1_127_reg_13928;
reg   [0:0] b1_127_reg_13928_pp0_iter1_reg;
wire   [0:0] b_93_fu_3100_p2;
reg   [0:0] b_93_reg_13933;
reg   [0:0] b_93_reg_13933_pp0_iter1_reg;
wire   [0:0] b0_37_fu_3208_p3;
reg   [0:0] b0_37_reg_13938;
reg   [0:0] b0_37_reg_13938_pp0_iter1_reg;
wire   [0:0] b0_33_fu_3278_p2;
reg   [0:0] b0_33_reg_13943;
reg   [0:0] b0_33_reg_13943_pp0_iter1_reg;
wire   [0:0] b1_129_fu_3284_p3;
reg   [0:0] b1_129_reg_13948;
reg   [0:0] b1_129_reg_13948_pp0_iter1_reg;
wire   [0:0] b_98_fu_3304_p2;
reg   [0:0] b_98_reg_13953;
reg   [0:0] b_98_reg_13953_pp0_iter1_reg;
wire   [0:0] b0_35_fu_3356_p3;
reg   [0:0] b0_35_reg_13958;
reg   [0:0] b0_35_reg_13958_pp0_iter1_reg;
wire   [0:0] b0_34_fu_3384_p2;
reg   [0:0] b0_34_reg_13963;
reg   [0:0] b0_34_reg_13963_pp0_iter1_reg;
wire   [0:0] b1_130_fu_3390_p3;
reg   [0:0] b1_130_reg_13968;
reg   [0:0] b1_130_reg_13968_pp0_iter1_reg;
wire   [0:0] b_102_fu_3410_p2;
reg   [0:0] b_102_reg_13973;
reg   [0:0] b_102_reg_13973_pp0_iter1_reg;
wire   [0:0] b1_131_fu_3456_p3;
reg   [0:0] b1_131_reg_13978;
reg   [0:0] b1_131_reg_13978_pp0_iter1_reg;
wire   [0:0] b_106_fu_3476_p2;
reg   [0:0] b_106_reg_13983;
reg   [0:0] b_106_reg_13983_pp0_iter1_reg;
wire   [0:0] b1_133_fu_3588_p3;
reg   [0:0] b1_133_reg_13988;
reg   [0:0] b1_133_reg_13988_pp0_iter1_reg;
wire   [0:0] b_111_fu_3608_p2;
reg   [0:0] b_111_reg_13993;
reg   [0:0] b_111_reg_13993_pp0_iter1_reg;
wire   [0:0] b0_39_fu_3660_p3;
reg   [0:0] b0_39_reg_13998;
reg   [0:0] b0_39_reg_13998_pp0_iter1_reg;
wire   [0:0] b0_38_fu_3688_p2;
reg   [0:0] b0_38_reg_14003;
reg   [0:0] b0_38_reg_14003_pp0_iter1_reg;
wire   [0:0] b1_134_fu_3694_p3;
reg   [0:0] b1_134_reg_14008;
reg   [0:0] b1_134_reg_14008_pp0_iter1_reg;
wire   [0:0] b_115_fu_3714_p2;
reg   [0:0] b_115_reg_14013;
reg   [0:0] b_115_reg_14013_pp0_iter1_reg;
wire   [0:0] b1_135_fu_3760_p3;
reg   [0:0] b1_135_reg_14018;
reg   [0:0] b1_135_reg_14018_pp0_iter1_reg;
wire   [0:0] b_119_fu_3780_p2;
reg   [0:0] b_119_reg_14023;
reg   [0:0] b_119_reg_14023_pp0_iter1_reg;
wire   [0:0] a0_329_fu_4156_p3;
reg   [0:0] a0_329_reg_14028;
reg   [0:0] a0_329_reg_14028_pp0_iter1_reg;
wire   [0:0] a1_307_fu_4164_p3;
reg   [0:0] a1_307_reg_14036;
reg   [0:0] a1_307_reg_14036_pp0_iter1_reg;
wire   [0:0] b_238_fu_4172_p2;
reg   [0:0] b_238_reg_14041;
reg   [0:0] b_238_reg_14041_pp0_iter1_reg;
wire   [0:0] a0_330_fu_4186_p3;
reg   [0:0] a0_330_reg_14046;
reg   [0:0] a0_330_reg_14046_pp0_iter1_reg;
wire   [0:0] a1_308_fu_4194_p3;
reg   [0:0] a1_308_reg_14052;
reg   [0:0] a1_308_reg_14052_pp0_iter1_reg;
wire   [0:0] a0_331_fu_4202_p2;
reg   [0:0] a0_331_reg_14057;
reg   [0:0] a0_331_reg_14057_pp0_iter1_reg;
wire   [0:0] a0_332_fu_4240_p3;
reg   [0:0] a0_332_reg_14062;
reg   [0:0] a0_332_reg_14062_pp0_iter1_reg;
wire   [0:0] a1_309_fu_4248_p3;
reg   [0:0] a1_309_reg_14069;
reg   [0:0] a1_309_reg_14069_pp0_iter1_reg;
wire   [0:0] b_264_fu_4256_p2;
reg   [0:0] b_264_reg_14074;
reg   [0:0] b_264_reg_14074_pp0_iter1_reg;
wire   [0:0] a0_333_fu_4270_p3;
reg   [0:0] a0_333_reg_14079;
reg   [0:0] a0_333_reg_14079_pp0_iter1_reg;
wire   [0:0] a1_310_fu_4278_p3;
reg   [0:0] a1_310_reg_14085;
reg   [0:0] a1_310_reg_14085_pp0_iter1_reg;
wire   [0:0] a0_334_fu_4286_p2;
reg   [0:0] a0_334_reg_14090;
reg   [0:0] a0_334_reg_14090_pp0_iter1_reg;
wire   [0:0] a1_311_fu_4354_p3;
reg   [0:0] a1_311_reg_14095;
reg   [0:0] a1_311_reg_14095_pp0_iter1_reg;
wire   [0:0] b_318_fu_4362_p2;
reg   [0:0] b_318_reg_14100;
reg   [0:0] b_318_reg_14100_pp0_iter1_reg;
wire   [0:0] a0_336_fu_4376_p3;
reg   [0:0] a0_336_reg_14105;
reg   [0:0] a0_336_reg_14105_pp0_iter1_reg;
wire   [0:0] a1_312_fu_4384_p3;
reg   [0:0] a1_312_reg_14111;
reg   [0:0] a1_312_reg_14111_pp0_iter1_reg;
wire   [0:0] a0_337_fu_4392_p2;
reg   [0:0] a0_337_reg_14116;
reg   [0:0] a0_337_reg_14116_pp0_iter1_reg;
wire   [0:0] a0_338_fu_4430_p3;
reg   [0:0] a0_338_reg_14121;
reg   [0:0] a0_338_reg_14121_pp0_iter1_reg;
wire   [0:0] a1_313_fu_4438_p3;
reg   [0:0] a1_313_reg_14128;
reg   [0:0] a1_313_reg_14128_pp0_iter1_reg;
wire   [0:0] b_344_fu_4446_p2;
reg   [0:0] b_344_reg_14133;
reg   [0:0] b_344_reg_14133_pp0_iter1_reg;
wire   [0:0] a0_343_fu_4756_p3;
reg   [0:0] a0_343_reg_14138;
reg   [0:0] a0_343_reg_14138_pp0_iter1_reg;
wire   [0:0] a1_318_fu_4764_p3;
reg   [0:0] a1_318_reg_14145;
reg   [0:0] a1_318_reg_14145_pp0_iter1_reg;
wire   [0:0] a0_361_fu_4772_p2;
reg   [0:0] a0_361_reg_14151;
reg   [0:0] a0_361_reg_14151_pp0_iter1_reg;
wire   [0:0] a0_360_fu_4816_p3;
reg   [0:0] a0_360_reg_14159;
reg   [0:0] a0_360_reg_14159_pp0_iter1_reg;
wire   [0:0] a0_346_fu_4922_p2;
reg   [0:0] a0_346_reg_14167;
reg   [0:0] a1_321_reg_14175;
wire   [0:0] b0_42_fu_5050_p2;
reg   [0:0] b0_42_reg_14181;
reg   [0:0] b0_42_reg_14181_pp0_iter1_reg;
reg   [0:0] b1_138_reg_14190;
reg   [0:0] b1_138_reg_14190_pp0_iter1_reg;
reg   [0:0] a0_348_reg_14197;
reg   [0:0] b0_44_reg_14204;
reg   [0:0] b0_44_reg_14204_pp0_iter1_reg;
reg   [0:0] a1_322_reg_14212;
reg   [0:0] b1_139_reg_14218;
reg   [0:0] b1_139_reg_14218_pp0_iter1_reg;
reg   [0:0] a1_323_reg_14225;
reg   [0:0] b1_140_reg_14231;
reg   [0:0] b1_140_reg_14231_pp0_iter1_reg;
reg   [0:0] a0_354_reg_14238;
reg   [0:0] b0_50_reg_14246;
reg   [0:0] b0_50_reg_14246_pp0_iter1_reg;
reg   [0:0] a1_325_reg_14255;
reg   [0:0] b1_142_reg_14261;
reg   [0:0] b1_142_reg_14261_pp0_iter1_reg;
reg   [0:0] a0_352_reg_14268;
reg   [0:0] b0_48_reg_14275;
reg   [0:0] b0_48_reg_14275_pp0_iter1_reg;
reg   [0:0] a1_326_reg_14283;
reg   [0:0] b1_143_reg_14289;
reg   [0:0] b1_143_reg_14289_pp0_iter1_reg;
reg   [0:0] a1_327_reg_14296;
reg   [0:0] b1_144_reg_14302;
reg   [0:0] b1_144_reg_14302_pp0_iter1_reg;
reg   [0:0] a1_329_reg_14309;
reg   [0:0] b1_146_reg_14315;
reg   [0:0] b1_146_reg_14315_pp0_iter1_reg;
reg   [0:0] a0_356_reg_14322;
reg   [0:0] b0_52_reg_14329;
reg   [0:0] b0_52_reg_14329_pp0_iter1_reg;
reg   [0:0] a1_330_reg_14337;
reg   [0:0] b1_147_reg_14343;
reg   [0:0] b1_147_reg_14343_pp0_iter1_reg;
reg   [0:0] a1_331_reg_14350;
reg   [0:0] b1_148_reg_14356;
reg   [0:0] b1_148_reg_14356_pp0_iter1_reg;
reg   [0:0] a0_357_reg_14363;
reg   [0:0] a0_357_reg_14363_pp0_iter1_reg;
reg   [0:0] a1_333_reg_14371;
reg   [0:0] a1_333_reg_14371_pp0_iter1_reg;
reg   [0:0] a0_358_reg_14378;
reg   [0:0] a0_358_reg_14378_pp0_iter1_reg;
reg   [0:0] a1_334_reg_14385;
reg   [0:0] a1_334_reg_14385_pp0_iter1_reg;
reg   [1:0] tmp_256_fu_5408_p4;
reg   [1:0] tmp_256_reg_14392;
reg   [0:0] a1_335_reg_14397;
reg   [0:0] a1_335_reg_14397_pp0_iter1_reg;
reg   [1:0] tmp_258_fu_5426_p4;
reg   [1:0] tmp_258_reg_14404;
reg   [0:0] b1_156_reg_14411;
reg   [0:0] b1_156_reg_14411_pp0_iter1_reg;
reg   [0:0] b1_158_reg_14417;
reg   [0:0] b1_158_reg_14417_pp0_iter1_reg;
reg   [0:0] b0_64_reg_14423;
reg   [0:0] b0_64_reg_14423_pp0_iter1_reg;
reg   [0:0] b1_159_reg_14430;
reg   [0:0] b1_159_reg_14430_pp0_iter1_reg;
reg   [0:0] b1_160_reg_14436;
reg   [0:0] b1_160_reg_14436_pp0_iter1_reg;
reg   [0:0] b1_161_reg_14442;
reg   [0:0] b1_161_reg_14442_pp0_iter1_reg;
reg   [0:0] b1_164_reg_14448;
reg   [0:0] b1_164_reg_14448_pp0_iter1_reg;
reg   [0:0] b1_166_reg_14454;
reg   [0:0] b1_166_reg_14454_pp0_iter1_reg;
reg   [0:0] b0_72_reg_14460;
reg   [0:0] b0_72_reg_14460_pp0_iter1_reg;
reg   [0:0] b1_167_reg_14467;
reg   [0:0] b1_167_reg_14467_pp0_iter1_reg;
reg   [0:0] b1_168_reg_14473;
reg   [0:0] b1_168_reg_14473_pp0_iter1_reg;
reg   [0:0] b1_170_reg_14479;
reg   [0:0] b1_170_reg_14479_pp0_iter1_reg;
reg   [0:0] b1_173_reg_14485;
reg   [0:0] b1_173_reg_14485_pp0_iter1_reg;
reg   [0:0] b0_79_reg_14491;
reg   [0:0] b0_79_reg_14491_pp0_iter1_reg;
reg   [0:0] b1_174_reg_14498;
reg   [0:0] b1_174_reg_14498_pp0_iter1_reg;
reg   [0:0] b1_175_reg_14504;
reg   [0:0] b1_175_reg_14504_pp0_iter1_reg;
reg   [0:0] b0_85_reg_14510;
reg   [0:0] b0_85_reg_14510_pp0_iter1_reg;
reg   [0:0] b1_177_reg_14518;
reg   [0:0] b1_177_reg_14518_pp0_iter1_reg;
reg   [0:0] b0_83_reg_14524;
reg   [0:0] b0_83_reg_14524_pp0_iter1_reg;
reg   [0:0] b1_178_reg_14531;
reg   [0:0] b1_178_reg_14531_pp0_iter1_reg;
reg   [0:0] b1_179_reg_14537;
reg   [0:0] b1_179_reg_14537_pp0_iter1_reg;
reg   [0:0] b1_181_reg_14543;
reg   [0:0] b1_181_reg_14543_pp0_iter1_reg;
reg   [0:0] b0_87_reg_14549;
reg   [0:0] b0_87_reg_14549_pp0_iter1_reg;
reg   [0:0] b1_182_reg_14556;
reg   [0:0] b1_182_reg_14556_pp0_iter1_reg;
reg   [0:0] b1_183_reg_14562;
reg   [0:0] b1_183_reg_14562_pp0_iter1_reg;
reg   [0:0] b1_185_reg_14568;
reg   [0:0] b1_185_reg_14568_pp0_iter1_reg;
reg   [0:0] b1_187_reg_14574;
reg   [0:0] b1_187_reg_14574_pp0_iter1_reg;
reg   [0:0] b0_93_reg_14580;
reg   [0:0] b0_93_reg_14580_pp0_iter1_reg;
reg   [0:0] b1_188_reg_14587;
reg   [0:0] b1_188_reg_14587_pp0_iter1_reg;
reg   [0:0] b1_189_reg_14593;
reg   [0:0] b1_189_reg_14593_pp0_iter1_reg;
reg   [0:0] b1_190_reg_14599;
reg   [0:0] b1_190_reg_14599_pp0_iter1_reg;
wire   [0:0] b_125_fu_5976_p2;
reg   [0:0] b_125_reg_14605;
wire   [0:0] b0_43_fu_6014_p2;
reg   [0:0] b0_43_reg_14610;
wire   [0:0] b_129_fu_6029_p2;
reg   [0:0] b_129_reg_14615;
wire   [0:0] b_133_fu_6072_p2;
reg   [0:0] b_133_reg_14620;
wire   [0:0] b0_46_fu_6156_p2;
reg   [0:0] b0_46_reg_14625;
wire   [0:0] b_138_fu_6171_p2;
reg   [0:0] b_138_reg_14630;
wire   [0:0] b0_47_fu_6211_p2;
reg   [0:0] b0_47_reg_14635;
wire   [0:0] b_142_fu_6227_p2;
reg   [0:0] b_142_reg_14640;
wire   [0:0] b_146_fu_6270_p2;
reg   [0:0] b_146_reg_14645;
wire   [0:0] b_151_fu_6358_p2;
reg   [0:0] b_151_reg_14650;
wire   [0:0] b0_51_fu_6396_p2;
reg   [0:0] b0_51_reg_14655;
wire   [0:0] b_155_fu_6411_p2;
reg   [0:0] b_155_reg_14660;
wire   [0:0] b_159_fu_6454_p2;
reg   [0:0] b_159_reg_14665;
wire   [0:0] b_198_fu_6624_p2;
reg   [0:0] b_198_reg_14670;
wire   [0:0] a0_359_fu_6635_p2;
reg   [0:0] a0_359_reg_14675;
wire   [0:0] b_224_fu_6659_p2;
reg   [0:0] b_224_reg_14680;
wire   [0:0] a0_364_fu_6769_p3;
reg   [0:0] a0_364_reg_14685;
wire   [0:0] a1_337_fu_6777_p3;
reg   [0:0] a1_337_reg_14691;
wire   [0:0] a0_370_fu_6785_p2;
reg   [0:0] a0_370_reg_14696;
wire   [0:0] b0_54_fu_6912_p2;
reg   [0:0] b0_54_reg_14701;
wire   [0:0] b1_150_fu_6918_p3;
reg   [0:0] b1_150_reg_14706;
wire   [0:0] b_164_fu_6938_p2;
reg   [0:0] b_164_reg_14711;
wire   [0:0] b0_56_fu_6990_p3;
reg   [0:0] b0_56_reg_14716;
wire   [0:0] b0_55_fu_7018_p2;
reg   [0:0] b0_55_reg_14721;
wire   [0:0] b1_151_fu_7024_p3;
reg   [0:0] b1_151_reg_14726;
wire   [0:0] b_168_fu_7044_p2;
reg   [0:0] b_168_reg_14731;
wire   [0:0] b1_152_fu_7090_p3;
reg   [0:0] b1_152_reg_14736;
wire   [0:0] b_172_fu_7110_p2;
reg   [0:0] b_172_reg_14741;
wire   [0:0] a0_369_fu_7206_p3;
reg   [0:0] a0_369_reg_14746;
wire   [0:0] a1_342_fu_7214_p3;
reg   [0:0] a1_342_reg_14752;
wire   [0:0] b_185_fu_7222_p2;
reg   [0:0] b_185_reg_14757;
wire   [0:0] a1_350_fu_7510_p2;
reg   [0:0] a1_350_reg_14762;
wire   [0:0] a0_379_fu_7516_p2;
reg   [0:0] a0_379_reg_14769;
wire   [0:0] a1_348_fu_7540_p2;
reg   [0:0] a1_348_reg_14777;
wire   [0:0] a0_377_fu_7546_p2;
reg   [0:0] a0_377_reg_14784;
wire   [0:0] a_233_fu_7552_p2;
reg   [0:0] a_233_reg_14792;
reg   [0:0] b1_154_reg_14798;
wire   [0:0] a_241_fu_7572_p2;
reg   [0:0] a_241_reg_14804;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_enable_reg_pp0_iter2;
wire    ap_block_pp0_stage0;
wire   [1:0] tmp_fu_266_p3;
wire   [1:0] a0_287_fu_224_p4;
wire   [1:0] xor_ln28_1_fu_274_p2;
wire   [1:0] a1_260_fu_234_p4;
wire   [3:0] tmp_1_fu_280_p3;
wire   [3:0] a0_286_fu_204_p4;
wire   [1:0] b0_88_fu_288_p4;
wire   [3:0] xor_ln28_2_fu_298_p2;
wire   [3:0] a1_259_fu_214_p4;
wire   [1:0] xor_ln28_23_fu_304_p2;
wire   [7:0] tmp_2_fu_310_p3;
wire   [7:0] a0_285_fu_184_p4;
wire   [5:0] tmp_95_fu_348_p3;
wire   [5:0] trunc_ln28_4_fu_338_p4;
wire   [1:0] b0_67_fu_328_p4;
wire   [3:0] b0_66_fu_318_p4;
wire   [7:0] xor_ln28_3_fu_356_p2;
wire   [7:0] a1_258_fu_194_p4;
wire   [3:0] xor_ln28_27_fu_382_p2;
wire   [1:0] xor_ln28_26_fu_376_p2;
wire   [5:0] xor_ln28_24_fu_370_p2;
wire   [15:0] tmp_3_fu_388_p3;
wire   [15:0] a0_284_fu_168_p1;
wire   [13:0] tmp_98_fu_432_p3;
wire   [13:0] trunc_ln68_1_fu_172_p1;
wire   [9:0] tmp_97_fu_424_p3;
wire   [9:0] trunc_ln68_2_fu_176_p1;
wire   [11:0] tmp_96_fu_416_p3;
wire   [11:0] trunc_ln68_3_fu_180_p1;
wire   [7:0] a0_289_fu_408_p1;
wire   [5:0] trunc_ln40_1_fu_474_p4;
wire   [5:0] trunc_ln70_4_fu_412_p1;
wire   [15:0] a0z1_fu_440_p2;
wire   [3:0] a0_290_fu_404_p1;
wire   [7:0] b0_fu_484_p2;
wire   [1:0] a0_291_fu_400_p1;
wire   [3:0] b0_1_fu_516_p2;
wire   [0:0] a0_292_fu_396_p1;
wire   [1:0] b0_2_fu_542_p2;
wire   [0:0] a1_265_fu_558_p3;
wire   [0:0] a_9_fu_586_p2;
wire   [0:0] z1_fu_598_p2;
wire   [0:0] z0_fu_580_p2;
wire   [0:0] z2_fu_604_p2;
wire   [0:0] xor_ln45_fu_610_p2;
wire   [0:0] xor_ln45_1_fu_616_p2;
wire   [1:0] a1_264_fu_532_p4;
wire   [1:0] b1_98_fu_548_p4;
wire   [0:0] a0_294_fu_630_p3;
wire   [1:0] a_11_fu_638_p2;
wire   [1:0] b_7_fu_652_p2;
wire   [0:0] a0_293_fu_658_p2;
wire   [0:0] a1_266_fu_664_p3;
wire   [0:0] a_13_fu_692_p2;
wire   [0:0] z1_1_fu_704_p2;
wire   [0:0] z0_2_fu_686_p2;
wire   [0:0] z2_1_fu_710_p2;
wire   [0:0] xor_ln45_2_fu_716_p2;
wire   [0:0] xor_ln45_3_fu_722_p2;
wire   [0:0] a1_267_fu_736_p3;
wire   [0:0] a_17_fu_758_p2;
wire   [0:0] z1_3_fu_770_p2;
wire   [0:0] z0_3_fu_752_p2;
wire   [0:0] z2_2_fu_776_p2;
wire   [0:0] a1_13_fu_782_p2;
wire   [0:0] a0_fu_788_p2;
wire   [0:0] xor_ln28_4_fu_802_p2;
wire   [1:0] z1_2_fu_728_p3;
wire   [1:0] z0_1_fu_622_p3;
wire   [1:0] z2_174_fu_794_p3;
wire   [1:0] tmp_7_fu_808_p3;
wire   [1:0] xor_ln45_7_fu_822_p2;
wire   [1:0] xor_ln45_6_fu_816_p2;
wire   [1:0] xor_ln45_8_fu_828_p2;
wire   [1:0] xor_ln45_9_fu_834_p2;
wire   [3:0] a1_263_fu_506_p4;
wire   [3:0] b1_97_fu_522_p4;
wire   [1:0] a0_299_fu_856_p4;
wire   [3:0] a_20_fu_866_p2;
wire   [1:0] b0_10_fu_880_p4;
wire   [3:0] b_15_fu_890_p2;
wire   [0:0] a0_300_fu_848_p3;
wire   [1:0] a0_295_fu_896_p2;
wire   [1:0] b0_6_fu_912_p2;
wire   [0:0] a0_296_fu_928_p2;
wire   [0:0] a1_269_fu_934_p3;
wire   [0:0] a_23_fu_962_p2;
wire   [0:0] z1_4_fu_974_p2;
wire   [0:0] z0_5_fu_956_p2;
wire   [0:0] z2_4_fu_980_p2;
wire   [0:0] xor_ln45_10_fu_986_p2;
wire   [0:0] xor_ln45_11_fu_992_p2;
wire   [1:0] a1_268_fu_902_p4;
wire   [1:0] b1_102_fu_918_p4;
wire   [0:0] a0_298_fu_1006_p3;
wire   [1:0] a_25_fu_1014_p2;
wire   [1:0] b_20_fu_1028_p2;
wire   [0:0] a0_297_fu_1034_p2;
wire   [0:0] a1_270_fu_1040_p3;
wire   [0:0] a_27_fu_1068_p2;
wire   [0:0] z1_5_fu_1080_p2;
wire   [0:0] z0_7_fu_1062_p2;
wire   [0:0] z2_5_fu_1086_p2;
wire   [0:0] xor_ln45_12_fu_1092_p2;
wire   [0:0] xor_ln45_13_fu_1098_p2;
wire   [0:0] a1_271_fu_1112_p3;
wire   [0:0] a_31_fu_1134_p2;
wire   [0:0] z1_7_fu_1146_p2;
wire   [0:0] z0_8_fu_1128_p2;
wire   [0:0] z2_6_fu_1152_p2;
wire   [0:0] a1_19_fu_1158_p2;
wire   [0:0] a0_16_fu_1164_p2;
wire   [0:0] xor_ln28_5_fu_1178_p2;
wire   [1:0] z1_6_fu_1104_p3;
wire   [1:0] z0_6_fu_998_p3;
wire   [1:0] z2_175_fu_1170_p3;
wire   [1:0] tmp_s_fu_1184_p3;
wire   [1:0] xor_ln45_17_fu_1198_p2;
wire   [1:0] xor_ln45_16_fu_1192_p2;
wire   [1:0] xor_ln45_18_fu_1204_p2;
wire   [1:0] xor_ln45_19_fu_1210_p2;
wire   [5:0] xor_ln40_1_fu_490_p2;
wire   [0:0] a1_273_fu_1244_p3;
wire   [0:0] a_37_fu_1266_p2;
wire   [0:0] z1_9_fu_1278_p2;
wire   [0:0] z0_9_fu_1260_p2;
wire   [0:0] z2_8_fu_1284_p2;
wire   [0:0] xor_ln45_20_fu_1290_p2;
wire   [0:0] xor_ln45_21_fu_1296_p2;
wire   [1:0] a1_272_fu_1224_p4;
wire   [1:0] b1_106_fu_1234_p4;
wire   [0:0] a0_302_fu_1310_p3;
wire   [1:0] a_39_fu_1318_p2;
wire   [1:0] b_33_fu_1332_p2;
wire   [0:0] a0_301_fu_1338_p2;
wire   [0:0] a1_274_fu_1344_p3;
wire   [0:0] a_41_fu_1372_p2;
wire   [0:0] z1_10_fu_1384_p2;
wire   [0:0] z0_11_fu_1366_p2;
wire   [0:0] z2_9_fu_1390_p2;
wire   [0:0] xor_ln45_22_fu_1396_p2;
wire   [0:0] xor_ln45_23_fu_1402_p2;
wire   [0:0] a1_275_fu_1416_p3;
wire   [0:0] a_45_fu_1438_p2;
wire   [0:0] z1_12_fu_1450_p2;
wire   [0:0] z0_12_fu_1432_p2;
wire   [0:0] z2_10_fu_1456_p2;
wire   [0:0] a1_24_fu_1462_p2;
wire   [0:0] a0_23_fu_1468_p2;
wire   [0:0] xor_ln28_6_fu_1482_p2;
wire   [1:0] z1_11_fu_1408_p3;
wire   [1:0] z0_10_fu_1302_p3;
wire   [1:0] z2_176_fu_1474_p3;
wire   [1:0] tmp_4_fu_1488_p3;
wire   [1:0] xor_ln45_27_fu_1502_p2;
wire   [1:0] xor_ln45_26_fu_1496_p2;
wire   [1:0] a1_276_fu_1508_p2;
wire   [1:0] a0_24_fu_1514_p2;
wire   [0:0] a0_25_fu_1528_p1;
wire   [0:0] a1_27_fu_1532_p3;
wire   [0:0] xor_ln28_7_fu_1540_p2;
wire   [1:0] tmp_5_fu_1546_p3;
wire   [1:0] xor_ln28_8_fu_1554_p2;
wire   [3:0] z1_8_fu_1216_p3;
wire   [3:0] z0_4_fu_840_p3;
wire   [3:0] z2_177_fu_1520_p3;
wire   [3:0] tmp_6_fu_1560_p3;
wire   [3:0] xor_ln45_31_fu_1574_p2;
wire   [3:0] xor_ln45_30_fu_1568_p2;
wire   [1:0] xor_ln45_39_fu_1586_p2;
wire   [1:0] xor_ln45_38_fu_1580_p2;
wire   [3:0] xor_ln45_32_fu_1592_p2;
wire   [3:0] xor_ln45_33_fu_1598_p2;
wire   [7:0] a1_262_fu_464_p4;
wire   [5:0] trunc_ln43_s_fu_1652_p4;
wire   [7:0] b1_fu_496_p4;
wire   [5:0] trunc_ln43_1_fu_1702_p4;
wire   [3:0] a0_316_fu_1642_p4;
wire   [7:0] a_50_fu_1662_p2;
wire   [3:0] b0_27_fu_1692_p4;
wire   [7:0] b_41_fu_1712_p2;
wire   [1:0] a0_317_fu_1632_p4;
wire   [3:0] a0_303_fu_1724_p2;
wire   [1:0] b0_28_fu_1682_p4;
wire   [3:0] b0_14_fu_1740_p2;
wire   [0:0] a0_318_fu_1624_p3;
wire   [1:0] a0_304_fu_1756_p2;
wire   [1:0] b0_15_fu_1772_p2;
wire   [0:0] a0_305_fu_1788_p2;
wire   [0:0] a1_279_fu_1794_p3;
wire   [0:0] a_54_fu_1822_p2;
wire   [0:0] z1_13_fu_1834_p2;
wire   [0:0] z0_14_fu_1816_p2;
wire   [0:0] z2_13_fu_1840_p2;
wire   [0:0] xor_ln45_34_fu_1846_p2;
wire   [0:0] xor_ln45_35_fu_1852_p2;
wire   [1:0] a1_278_fu_1762_p4;
wire   [1:0] b1_111_fu_1778_p4;
wire   [0:0] a0_307_fu_1866_p3;
wire   [1:0] a_56_fu_1874_p2;
wire   [1:0] b_47_fu_1888_p2;
wire   [0:0] a0_306_fu_1894_p2;
wire   [0:0] a1_280_fu_1900_p3;
wire   [0:0] a_58_fu_1928_p2;
wire   [0:0] z1_14_fu_1940_p2;
wire   [0:0] z0_16_fu_1922_p2;
wire   [0:0] z2_14_fu_1946_p2;
wire   [0:0] xor_ln45_36_fu_1952_p2;
wire   [0:0] xor_ln45_37_fu_1958_p2;
wire   [0:0] a1_281_fu_1972_p3;
wire   [0:0] a_62_fu_1994_p2;
wire   [0:0] z1_16_fu_2006_p2;
wire   [0:0] z0_17_fu_1988_p2;
wire   [0:0] z2_15_fu_2012_p2;
wire   [0:0] a1_34_fu_2018_p2;
wire   [0:0] a0_36_fu_2024_p2;
wire   [0:0] xor_ln28_9_fu_2038_p2;
wire   [1:0] z1_15_fu_1964_p3;
wire   [1:0] z0_15_fu_1858_p3;
wire   [1:0] z2_178_fu_2030_p3;
wire   [1:0] tmp_8_fu_2044_p3;
wire   [1:0] xor_ln45_51_fu_2058_p2;
wire   [1:0] xor_ln45_50_fu_2052_p2;
wire   [1:0] xor_ln45_42_fu_2064_p2;
wire   [1:0] xor_ln45_43_fu_2070_p2;
wire   [3:0] a1_277_fu_1730_p4;
wire   [3:0] b1_110_fu_1746_p4;
wire   [1:0] a0_312_fu_2092_p4;
wire   [3:0] a_65_fu_2102_p2;
wire   [1:0] b0_23_fu_2116_p4;
wire   [3:0] b_55_fu_2126_p2;
wire   [0:0] a0_313_fu_2084_p3;
wire   [1:0] a0_308_fu_2132_p2;
wire   [1:0] b0_19_fu_2148_p2;
wire   [0:0] a0_309_fu_2164_p2;
wire   [0:0] a1_283_fu_2170_p3;
wire   [0:0] a_68_fu_2198_p2;
wire   [0:0] z1_17_fu_2210_p2;
wire   [0:0] z0_19_fu_2192_p2;
wire   [0:0] z2_17_fu_2216_p2;
wire   [0:0] xor_ln45_44_fu_2222_p2;
wire   [0:0] xor_ln45_45_fu_2228_p2;
wire   [1:0] a1_282_fu_2138_p4;
wire   [1:0] b1_115_fu_2154_p4;
wire   [0:0] a0_311_fu_2242_p3;
wire   [1:0] a_70_fu_2250_p2;
wire   [1:0] b_60_fu_2264_p2;
wire   [0:0] a0_310_fu_2270_p2;
wire   [0:0] a1_284_fu_2276_p3;
wire   [0:0] a_72_fu_2304_p2;
wire   [0:0] z1_18_fu_2316_p2;
wire   [0:0] z0_21_fu_2298_p2;
wire   [0:0] z2_18_fu_2322_p2;
wire   [0:0] xor_ln45_46_fu_2328_p2;
wire   [0:0] xor_ln45_47_fu_2334_p2;
wire   [0:0] a1_285_fu_2348_p3;
wire   [0:0] a_76_fu_2370_p2;
wire   [0:0] z1_20_fu_2382_p2;
wire   [0:0] z0_22_fu_2364_p2;
wire   [0:0] z2_19_fu_2388_p2;
wire   [0:0] a1_40_fu_2394_p2;
wire   [0:0] a0_45_fu_2400_p2;
wire   [0:0] xor_ln28_10_fu_2414_p2;
wire   [1:0] z1_19_fu_2340_p3;
wire   [1:0] z0_20_fu_2234_p3;
wire   [1:0] z2_179_fu_2406_p3;
wire   [1:0] tmp_9_fu_2420_p3;
wire   [1:0] xor_ln45_61_fu_2434_p2;
wire   [1:0] xor_ln45_60_fu_2428_p2;
wire   [1:0] xor_ln45_52_fu_2440_p2;
wire   [1:0] xor_ln45_53_fu_2446_p2;
wire   [5:0] xor_ln43_14_fu_1668_p2;
wire   [5:0] xor_ln33_fu_1718_p2;
wire   [0:0] a1_287_fu_2480_p3;
wire   [0:0] a_82_fu_2502_p2;
wire   [0:0] z1_22_fu_2514_p2;
wire   [0:0] z0_23_fu_2496_p2;
wire   [0:0] z2_21_fu_2520_p2;
wire   [0:0] xor_ln45_54_fu_2526_p2;
wire   [0:0] xor_ln45_55_fu_2532_p2;
wire   [1:0] a1_286_fu_2460_p4;
wire   [1:0] b1_119_fu_2470_p4;
wire   [0:0] a0_315_fu_2546_p3;
wire   [1:0] a_84_fu_2554_p2;
wire   [1:0] b_73_fu_2568_p2;
wire   [0:0] a0_314_fu_2574_p2;
wire   [0:0] a1_288_fu_2580_p3;
wire   [0:0] a_86_fu_2608_p2;
wire   [0:0] z1_23_fu_2620_p2;
wire   [0:0] z0_25_fu_2602_p2;
wire   [0:0] z2_22_fu_2626_p2;
wire   [0:0] xor_ln45_56_fu_2632_p2;
wire   [0:0] xor_ln45_57_fu_2638_p2;
wire   [0:0] a1_289_fu_2652_p3;
wire   [0:0] a_90_fu_2674_p2;
wire   [0:0] z1_25_fu_2686_p2;
wire   [0:0] z0_26_fu_2668_p2;
wire   [0:0] z2_23_fu_2692_p2;
wire   [0:0] a1_46_fu_2698_p2;
wire   [0:0] a0_49_fu_2704_p2;
wire   [0:0] xor_ln28_11_fu_2718_p2;
wire   [1:0] z1_24_fu_2644_p3;
wire   [1:0] z0_24_fu_2538_p3;
wire   [1:0] z2_180_fu_2710_p3;
wire   [1:0] tmp_10_fu_2724_p3;
wire   [1:0] xor_ln45_65_fu_2738_p2;
wire   [1:0] xor_ln45_64_fu_2732_p2;
wire   [1:0] a1_290_fu_2744_p2;
wire   [1:0] a0_50_fu_2750_p2;
wire   [0:0] a0_52_fu_2764_p1;
wire   [0:0] a1_49_fu_2768_p3;
wire   [0:0] xor_ln28_12_fu_2776_p2;
wire   [1:0] tmp_11_fu_2782_p3;
wire   [1:0] xor_ln28_13_fu_2790_p2;
wire   [3:0] z1_21_fu_2452_p3;
wire   [3:0] z0_18_fu_2076_p3;
wire   [3:0] z2_181_fu_2756_p3;
wire   [3:0] tmp_12_fu_2796_p3;
wire   [3:0] xor_ln45_75_fu_2810_p2;
wire   [3:0] xor_ln45_74_fu_2804_p2;
wire   [1:0] xor_ln45_83_fu_2822_p2;
wire   [1:0] xor_ln45_82_fu_2816_p2;
wire   [3:0] xor_ln45_66_fu_2828_p2;
wire   [3:0] xor_ln45_67_fu_2834_p2;
wire   [11:0] xor_ln70_3_fu_458_p2;
wire   [9:0] xor_ln70_2_fu_452_p2;
wire   [0:0] a1_293_fu_2900_p3;
wire   [0:0] a_99_fu_2922_p2;
wire   [0:0] z1_27_fu_2934_p2;
wire   [0:0] z0_27_fu_2916_p2;
wire   [0:0] z2_26_fu_2940_p2;
wire   [0:0] xor_ln45_68_fu_2946_p2;
wire   [0:0] xor_ln45_69_fu_2952_p2;
wire   [1:0] a1_292_fu_2880_p4;
wire   [1:0] b1_124_fu_2890_p4;
wire   [0:0] a0_320_fu_2966_p3;
wire   [1:0] a_101_fu_2974_p2;
wire   [1:0] b_87_fu_2988_p2;
wire   [0:0] a0_319_fu_2994_p2;
wire   [0:0] a1_294_fu_3000_p3;
wire   [0:0] a_103_fu_3028_p2;
wire   [0:0] z1_28_fu_3040_p2;
wire   [0:0] z0_29_fu_3022_p2;
wire   [0:0] z2_27_fu_3046_p2;
wire   [0:0] xor_ln45_70_fu_3052_p2;
wire   [0:0] xor_ln45_71_fu_3058_p2;
wire   [0:0] a1_295_fu_3072_p3;
wire   [0:0] a_107_fu_3094_p2;
wire   [0:0] z1_30_fu_3106_p2;
wire   [0:0] z0_30_fu_3088_p2;
wire   [0:0] z2_28_fu_3112_p2;
wire   [0:0] a1_56_fu_3118_p2;
wire   [0:0] a0_57_fu_3124_p2;
wire   [0:0] xor_ln28_14_fu_3138_p2;
wire   [1:0] z1_29_fu_3064_p3;
wire   [1:0] z0_28_fu_2958_p3;
wire   [1:0] z2_182_fu_3130_p3;
wire   [1:0] tmp_13_fu_3144_p3;
wire   [1:0] xor_ln45_95_fu_3158_p2;
wire   [1:0] xor_ln45_94_fu_3152_p2;
wire   [1:0] xor_ln45_76_fu_3164_p2;
wire   [1:0] xor_ln45_77_fu_3170_p2;
wire   [3:0] a1_291_fu_2860_p4;
wire   [3:0] b1_123_fu_2870_p4;
wire   [1:0] a0_325_fu_3192_p4;
wire   [3:0] a_110_fu_3202_p2;
wire   [1:0] b0_36_fu_3216_p4;
wire   [3:0] b_95_fu_3226_p2;
wire   [0:0] a0_326_fu_3184_p3;
wire   [1:0] a0_321_fu_3232_p2;
wire   [1:0] b0_32_fu_3248_p2;
wire   [0:0] a0_322_fu_3264_p2;
wire   [0:0] a1_297_fu_3270_p3;
wire   [0:0] a_113_fu_3298_p2;
wire   [0:0] z1_31_fu_3310_p2;
wire   [0:0] z0_32_fu_3292_p2;
wire   [0:0] z2_30_fu_3316_p2;
wire   [0:0] xor_ln45_78_fu_3322_p2;
wire   [0:0] xor_ln45_79_fu_3328_p2;
wire   [1:0] a1_296_fu_3238_p4;
wire   [1:0] b1_128_fu_3254_p4;
wire   [0:0] a0_324_fu_3342_p3;
wire   [1:0] a_115_fu_3350_p2;
wire   [1:0] b_100_fu_3364_p2;
wire   [0:0] a0_323_fu_3370_p2;
wire   [0:0] a1_298_fu_3376_p3;
wire   [0:0] a_117_fu_3404_p2;
wire   [0:0] z1_32_fu_3416_p2;
wire   [0:0] z0_34_fu_3398_p2;
wire   [0:0] z2_31_fu_3422_p2;
wire   [0:0] xor_ln45_80_fu_3428_p2;
wire   [0:0] xor_ln45_81_fu_3434_p2;
wire   [0:0] a1_299_fu_3448_p3;
wire   [0:0] a_121_fu_3470_p2;
wire   [0:0] z1_34_fu_3482_p2;
wire   [0:0] z0_35_fu_3464_p2;
wire   [0:0] z2_32_fu_3488_p2;
wire   [0:0] a1_61_fu_3494_p2;
wire   [0:0] a0_64_fu_3500_p2;
wire   [0:0] xor_ln28_15_fu_3514_p2;
wire   [1:0] z1_33_fu_3440_p3;
wire   [1:0] z0_33_fu_3334_p3;
wire   [1:0] z2_183_fu_3506_p3;
wire   [1:0] tmp_14_fu_3520_p3;
wire   [1:0] xor_ln45_99_fu_3534_p2;
wire   [1:0] xor_ln45_98_fu_3528_p2;
wire   [1:0] xor_ln45_86_fu_3540_p2;
wire   [1:0] xor_ln45_87_fu_3546_p2;
wire   [13:0] xor_ln70_1_fu_446_p2;
wire   [0:0] a1_301_fu_3580_p3;
wire   [0:0] a_127_fu_3602_p2;
wire   [0:0] z1_36_fu_3614_p2;
wire   [0:0] z0_36_fu_3596_p2;
wire   [0:0] z2_34_fu_3620_p2;
wire   [0:0] xor_ln45_88_fu_3626_p2;
wire   [0:0] xor_ln45_89_fu_3632_p2;
wire   [1:0] a1_300_fu_3560_p4;
wire   [1:0] b1_132_fu_3570_p4;
wire   [0:0] a0_328_fu_3646_p3;
wire   [1:0] a_129_fu_3654_p2;
wire   [1:0] b_113_fu_3668_p2;
wire   [0:0] a0_327_fu_3674_p2;
wire   [0:0] a1_302_fu_3680_p3;
wire   [0:0] a_131_fu_3708_p2;
wire   [0:0] z1_37_fu_3720_p2;
wire   [0:0] z0_38_fu_3702_p2;
wire   [0:0] z2_35_fu_3726_p2;
wire   [0:0] xor_ln45_90_fu_3732_p2;
wire   [0:0] xor_ln45_91_fu_3738_p2;
wire   [0:0] a1_303_fu_3752_p3;
wire   [0:0] a_135_fu_3774_p2;
wire   [0:0] z1_39_fu_3786_p2;
wire   [0:0] z0_39_fu_3768_p2;
wire   [0:0] z2_36_fu_3792_p2;
wire   [0:0] a1_66_fu_3798_p2;
wire   [0:0] a0_69_fu_3804_p2;
wire   [0:0] xor_ln28_16_fu_3818_p2;
wire   [1:0] z1_38_fu_3744_p3;
wire   [1:0] z0_37_fu_3638_p3;
wire   [1:0] z2_184_fu_3810_p3;
wire   [1:0] tmp_15_fu_3824_p3;
wire   [1:0] xor_ln45_103_fu_3838_p2;
wire   [1:0] xor_ln45_102_fu_3832_p2;
wire   [1:0] a1_304_fu_3844_p2;
wire   [1:0] a0_70_fu_3850_p2;
wire   [0:0] a0_72_fu_3864_p1;
wire   [0:0] a1_68_fu_3868_p3;
wire   [0:0] xor_ln28_17_fu_3876_p2;
wire   [1:0] tmp_16_fu_3882_p3;
wire   [1:0] xor_ln28_18_fu_3890_p2;
wire   [3:0] z1_35_fu_3552_p3;
wire   [3:0] z0_31_fu_3176_p3;
wire   [3:0] z2_185_fu_3856_p3;
wire   [3:0] tmp_17_fu_3896_p3;
wire   [3:0] xor_ln45_113_fu_3910_p2;
wire   [3:0] xor_ln45_112_fu_3904_p2;
wire   [1:0] xor_ln45_121_fu_3922_p2;
wire   [1:0] xor_ln45_120_fu_3916_p2;
wire   [3:0] a1_305_fu_3928_p2;
wire   [3:0] a0_73_fu_3934_p2;
wire   [0:0] a0_76_fu_3974_p3;
wire   [0:0] a1_71_fu_3982_p3;
wire   [0:0] xor_ln28_19_fu_3990_p2;
wire   [1:0] a0_74_fu_3960_p1;
wire   [1:0] tmp_18_fu_3996_p3;
wire   [1:0] xor_ln28_20_fu_4004_p2;
wire   [1:0] a1_306_fu_3964_p4;
wire   [3:0] tmp_19_fu_4010_p3;
wire   [1:0] xor_ln45_131_fu_3946_p2;
wire   [3:0] xor_ln28_21_fu_4018_p2;
wire   [1:0] xor_ln45_40_fu_1604_p2;
wire   [1:0] xor_ln45_85_fu_2846_p2;
wire   [7:0] z1_26_fu_2852_p3;
wire   [7:0] z0_13_fu_1616_p3;
wire   [1:0] xor_ln28_28_fu_4024_p2;
wire   [1:0] xor_ln45_130_fu_3940_p2;
wire   [7:0] z2_186_fu_3952_p3;
wire   [7:0] tmp_20_fu_4030_p3;
wire   [1:0] xor_ln45_84_fu_2840_p2;
wire   [1:0] xor_ln45_41_fu_1610_p2;
wire   [5:0] tmp_100_fu_4046_p3;
wire   [5:0] tmp_99_fu_4038_p3;
wire   [5:0] tmp_102_fu_4068_p3;
wire   [5:0] tmp_101_fu_4060_p3;
wire   [7:0] xor_ln45_133_fu_4076_p2;
wire   [7:0] xor_ln45_132_fu_4054_p2;
wire   [5:0] xor_ln45_145_fu_4112_p2;
wire   [5:0] xor_ln45_144_fu_4106_p2;
wire   [1:0] xor_ln45_137_fu_4100_p2;
wire   [1:0] xor_ln45_136_fu_4094_p2;
wire   [3:0] xor_ln45_135_fu_4088_p2;
wire   [3:0] xor_ln45_134_fu_4082_p2;
wire   [7:0] xor_ln45_104_fu_4118_p2;
wire   [7:0] xor_ln45_105_fu_4124_p2;
wire   [1:0] a1_sqr_fu_4208_p3;
wire   [1:0] a0_sqr_1_fu_4178_p3;
reg   [1:0] tmp_208_fu_4222_p4;
wire   [1:0] xor_ln59_2_fu_4216_p2;
wire   [1:0] a1_sqr_25_fu_4292_p3;
wire   [1:0] a0_sqr_5_fu_4262_p3;
reg   [1:0] tmp_213_fu_4306_p4;
wire   [1:0] a0_86_fu_4300_p2;
wire   [1:0] tmp_22_fu_4324_p3;
wire   [3:0] a1_sqr_26_fu_4316_p3;
wire   [3:0] a0_sqr_3_fu_4232_p3;
wire   [1:0] xor_ln28_25_fu_4332_p2;
wire   [3:0] xor_ln59_6_fu_4338_p2;
wire   [1:0] a1_sqr_27_fu_4398_p3;
wire   [1:0] a0_sqr_9_fu_4368_p3;
reg   [1:0] tmp_217_fu_4412_p4;
wire   [1:0] xor_ln59_9_fu_4406_p2;
wire   [1:0] a1_sqr_28_fu_4460_p3;
wire   [1:0] a0_sqr_13_fu_4452_p3;
reg   [1:0] a1_314_fu_4474_p4;
wire   [1:0] a0_94_fu_4468_p2;
wire   [1:0] tmp_23_fu_4492_p3;
wire   [3:0] a1_sqr_29_fu_4484_p3;
wire   [3:0] a0_sqr_11_fu_4422_p3;
wire   [1:0] a1_315_fu_4500_p2;
wire   [3:0] a0_96_fu_4506_p2;
wire   [0:0] a0_98_fu_4522_p1;
wire   [0:0] a1_88_fu_4526_p3;
wire   [0:0] xor_ln28_30_fu_4534_p2;
wire   [1:0] tmp_24_fu_4540_p3;
wire   [1:0] xor_ln28_31_fu_4548_p2;
wire   [3:0] tmp_25_fu_4554_p3;
wire   [7:0] a1_sqr_30_fu_4512_p4;
wire   [7:0] a0_sqr_7_fu_4344_p4;
wire   [3:0] xor_ln28_32_fu_4568_p2;
wire   [7:0] xor_ln59_13_fu_4590_p2;
wire   [3:0] xor_ln45_152_fu_4142_p2;
wire   [1:0] xor_ln45_147_fu_4136_p2;
wire   [5:0] xor_ln45_146_fu_4130_p2;
wire   [1:0] xor_ln59_14_fu_4596_p2;
wire   [15:0] tmp_26_fu_4602_p5;
wire   [15:0] tmp_21_fu_4148_p3;
wire   [13:0] tmp_110_fu_4656_p5;
wire   [13:0] tmp_109_fu_4648_p3;
wire   [9:0] tmp_108_fu_4640_p3;
wire   [9:0] tmp_107_fu_4632_p3;
wire   [11:0] tmp_106_fu_4622_p4;
wire   [11:0] tmp_105_fu_4614_p3;
wire   [5:0] tmp_104_fu_4582_p3;
wire   [5:0] tmp_103_fu_4574_p3;
wire   [5:0] xor_ln68_1_fu_4698_p2;
wire   [5:0] xor_ln68_fu_4692_p2;
wire   [11:0] xor_ln71_3_fu_4686_p2;
wire   [15:0] delta_fu_4668_p2;
wire   [1:0] a0_342_fu_4736_p4;
wire   [1:0] tmp_27_fu_4778_p3;
wire   [1:0] xor_ln28_34_fu_4786_p2;
wire   [1:0] a1_317_fu_4746_p4;
wire   [3:0] a0_341_fu_4716_p4;
wire   [3:0] tmp_28_fu_4792_p3;
wire   [1:0] b0_59_fu_4800_p4;
wire   [3:0] xor_ln28_35_fu_4810_p2;
wire   [3:0] a1_316_fu_4726_p4;
wire   [0:0] xor_ln70_4_fu_4844_p2;
wire   [0:0] xor_ln70_fu_4838_p2;
wire   [0:0] xor_ln70_7_fu_4862_p2;
wire   [0:0] xor_ln70_6_fu_4856_p2;
wire   [0:0] xor_ln70_8_fu_4868_p2;
wire   [0:0] xor_ln70_5_fu_4850_p2;
wire   [0:0] xor_ln70_11_fu_4886_p2;
wire   [0:0] xor_ln70_10_fu_4880_p2;
wire   [0:0] xor_ln70_14_fu_4904_p2;
wire   [0:0] xor_ln70_13_fu_4898_p2;
wire   [0:0] xor_ln70_15_fu_4910_p2;
wire   [0:0] xor_ln70_12_fu_4892_p2;
wire   [0:0] xor_ln70_16_fu_4916_p2;
wire   [0:0] xor_ln70_9_fu_4874_p2;
wire   [1:0] xor_ln28_33_fu_4562_p2;
wire   [1:0] xor_ln70_18_fu_4928_p2;
wire   [1:0] xor_ln70_21_fu_4940_p2;
wire   [1:0] xor_ln70_20_fu_4934_p2;
wire   [3:0] xor_ln70_24_fu_4958_p2;
wire   [3:0] xor_ln70_23_fu_4952_p2;
wire   [1:0] xor_ln28_42_fu_4824_p2;
wire   [7:0] tmp_29_fu_4830_p3;
wire   [7:0] a0_340_fu_4704_p2;
wire   [5:0] tmp_111_fu_4970_p3;
wire   [5:0] xor_ln68_3_fu_4710_p2;
wire   [3:0] a0_344_fu_4964_p2;
wire   [7:0] a0z1_1_fu_4978_p2;
wire   [1:0] a0_345_fu_4946_p2;
wire   [3:0] b0_40_fu_5000_p2;
wire   [1:0] b0_41_fu_5026_p2;
wire   [1:0] a1_320_fu_5016_p4;
wire   [1:0] b1_137_fu_5032_p4;
wire   [1:0] a_161_fu_5072_p2;
wire   [1:0] b_127_fu_5086_p2;
wire   [3:0] a1_319_fu_4990_p4;
wire   [3:0] b1_136_fu_5006_p4;
wire   [1:0] a0_353_fu_5132_p4;
wire   [3:0] a_170_fu_5142_p2;
wire   [1:0] b0_49_fu_5156_p4;
wire   [3:0] b_135_fu_5166_p2;
wire   [1:0] a0_349_fu_5172_p2;
wire   [1:0] b0_45_fu_5188_p2;
wire   [1:0] a1_324_fu_5178_p4;
wire   [1:0] b1_141_fu_5194_p4;
wire   [1:0] a_175_fu_5228_p2;
wire   [1:0] b_140_fu_5242_p2;
wire   [5:0] xor_ln70_27_fu_4984_p2;
wire   [1:0] a1_328_fu_5280_p4;
wire   [1:0] b1_145_fu_5290_p4;
wire   [1:0] a_189_fu_5324_p2;
wire   [1:0] b_153_fu_5338_p2;
wire   [9:0] xor_ln71_2_fu_4680_p2;
wire   [13:0] xor_ln71_1_fu_4674_p2;
wire   [1:0] b1_155_fu_5436_p4;
wire   [1:0] b_200_fu_5446_p2;
wire   [3:0] b_208_fu_5460_p2;
wire   [1:0] b0_61_fu_5466_p2;
wire   [1:0] b1_157_fu_5472_p4;
wire   [1:0] b_213_fu_5498_p2;
wire   [1:0] b_226_fu_5520_p2;
wire   [1:0] b1_163_fu_5544_p4;
wire   [1:0] b_240_fu_5554_p2;
wire   [3:0] b1_162_fu_5534_p4;
wire   [1:0] b0_73_fu_5568_p4;
wire   [3:0] b_248_fu_5578_p2;
wire   [1:0] b0_69_fu_5584_p2;
wire   [1:0] b1_165_fu_5590_p4;
wire   [1:0] b_253_fu_5616_p2;
wire   [1:0] b1_169_fu_5638_p4;
wire   [1:0] b_266_fu_5648_p2;
wire   [7:0] b_274_fu_5662_p2;
wire   [3:0] b0_75_fu_5674_p2;
wire   [1:0] b0_76_fu_5690_p2;
wire   [1:0] b1_172_fu_5696_p4;
wire   [1:0] b_280_fu_5722_p2;
wire   [3:0] b1_171_fu_5680_p4;
wire   [1:0] b0_84_fu_5752_p4;
wire   [3:0] b_288_fu_5762_p2;
wire   [1:0] b0_80_fu_5768_p2;
wire   [1:0] b1_176_fu_5774_p4;
wire   [1:0] b_293_fu_5800_p2;
wire   [5:0] xor_ln33_1_fu_5668_p2;
wire   [1:0] b1_180_fu_5822_p4;
wire   [1:0] b_306_fu_5848_p2;
wire   [1:0] b1_184_fu_5870_p4;
wire   [1:0] b_320_fu_5880_p2;
wire   [3:0] b_328_fu_5894_p2;
wire   [1:0] b0_90_fu_5900_p2;
wire   [1:0] b1_186_fu_5906_p4;
wire   [1:0] b_333_fu_5932_p2;
wire   [1:0] b_346_fu_5954_p2;
wire   [0:0] a_159_fu_5972_p2;
wire   [0:0] z1_40_fu_5980_p2;
wire   [0:0] z0_40_fu_5968_p2;
wire   [0:0] z2_40_fu_5986_p2;
wire   [0:0] xor_ln45_106_fu_5990_p2;
wire   [0:0] xor_ln45_107_fu_5996_p2;
wire   [0:0] a0_347_fu_6010_p2;
wire   [0:0] a_163_fu_6024_p2;
wire   [0:0] z1_41_fu_6034_p2;
wire   [0:0] z0_42_fu_6018_p2;
wire   [0:0] z2_41_fu_6040_p2;
wire   [0:0] xor_ln45_108_fu_6044_p2;
wire   [0:0] xor_ln45_109_fu_6050_p2;
wire   [0:0] a_167_fu_6068_p2;
wire   [0:0] z1_43_fu_6076_p2;
wire   [0:0] z0_43_fu_6064_p2;
wire   [0:0] z2_42_fu_6082_p2;
wire   [0:0] a1_98_fu_6086_p2;
wire   [0:0] a0_111_fu_6092_p2;
wire   [0:0] xor_ln28_36_fu_6106_p2;
wire   [1:0] z1_42_fu_6056_p3;
wire   [1:0] z0_41_fu_6002_p3;
wire   [1:0] z2_187_fu_6098_p3;
wire   [1:0] tmp_30_fu_6112_p3;
wire   [1:0] xor_ln45_160_fu_6126_p2;
wire   [1:0] xor_ln45_155_fu_6120_p2;
wire   [1:0] xor_ln45_114_fu_6132_p2;
wire   [1:0] xor_ln45_115_fu_6138_p2;
wire   [0:0] a0_350_fu_6152_p2;
wire   [0:0] a_173_fu_6166_p2;
wire   [0:0] z1_44_fu_6176_p2;
wire   [0:0] z0_45_fu_6160_p2;
wire   [0:0] z2_44_fu_6182_p2;
wire   [0:0] xor_ln45_116_fu_6186_p2;
wire   [0:0] xor_ln45_117_fu_6192_p2;
wire   [0:0] a0_351_fu_6206_p2;
wire   [0:0] a_177_fu_6222_p2;
wire   [0:0] z1_45_fu_6232_p2;
wire   [0:0] z0_47_fu_6216_p2;
wire   [0:0] z2_45_fu_6238_p2;
wire   [0:0] xor_ln45_118_fu_6242_p2;
wire   [0:0] xor_ln45_119_fu_6248_p2;
wire   [0:0] a_181_fu_6266_p2;
wire   [0:0] z1_47_fu_6274_p2;
wire   [0:0] z0_48_fu_6262_p2;
wire   [0:0] z2_46_fu_6280_p2;
wire   [0:0] a1_103_fu_6284_p2;
wire   [0:0] a0_117_fu_6290_p2;
wire   [0:0] xor_ln28_37_fu_6304_p2;
wire   [1:0] z1_46_fu_6254_p3;
wire   [1:0] z0_46_fu_6198_p3;
wire   [1:0] z2_188_fu_6296_p3;
wire   [1:0] tmp_31_fu_6310_p3;
wire   [1:0] xor_ln45_164_fu_6324_p2;
wire   [1:0] xor_ln45_163_fu_6318_p2;
wire   [1:0] xor_ln45_124_fu_6330_p2;
wire   [1:0] xor_ln45_125_fu_6336_p2;
wire   [0:0] a_187_fu_6354_p2;
wire   [0:0] z1_49_fu_6362_p2;
wire   [0:0] z0_49_fu_6350_p2;
wire   [0:0] z2_48_fu_6368_p2;
wire   [0:0] xor_ln45_126_fu_6372_p2;
wire   [0:0] xor_ln45_127_fu_6378_p2;
wire   [0:0] a0_355_fu_6392_p2;
wire   [0:0] a_191_fu_6406_p2;
wire   [0:0] z1_50_fu_6416_p2;
wire   [0:0] z0_51_fu_6400_p2;
wire   [0:0] z2_49_fu_6422_p2;
wire   [0:0] xor_ln45_128_fu_6426_p2;
wire   [0:0] xor_ln45_129_fu_6432_p2;
wire   [0:0] a_195_fu_6450_p2;
wire   [0:0] z1_52_fu_6458_p2;
wire   [0:0] z0_52_fu_6446_p2;
wire   [0:0] z2_50_fu_6464_p2;
wire   [0:0] a1_109_fu_6468_p2;
wire   [0:0] a0_128_fu_6474_p2;
wire   [0:0] xor_ln28_38_fu_6488_p2;
wire   [1:0] z1_51_fu_6438_p3;
wire   [1:0] z0_50_fu_6384_p3;
wire   [1:0] z2_189_fu_6480_p3;
wire   [1:0] tmp_32_fu_6494_p3;
wire   [1:0] xor_ln45_172_fu_6508_p2;
wire   [1:0] xor_ln45_171_fu_6502_p2;
wire   [1:0] a1_332_fu_6514_p2;
wire   [1:0] a0_129_fu_6520_p2;
wire   [0:0] a0_130_fu_6534_p1;
wire   [0:0] a1_111_fu_6538_p3;
wire   [0:0] xor_ln28_39_fu_6546_p2;
wire   [1:0] tmp_33_fu_6552_p3;
wire   [1:0] xor_ln28_40_fu_6560_p2;
wire   [3:0] z1_48_fu_6342_p3;
wire   [3:0] z0_44_fu_6144_p3;
wire   [3:0] z2_190_fu_6526_p3;
wire   [3:0] tmp_34_fu_6566_p3;
wire   [3:0] xor_ln45_180_fu_6580_p2;
wire   [3:0] xor_ln45_175_fu_6574_p2;
wire   [1:0] xor_ln45_182_fu_6592_p2;
wire   [1:0] xor_ln45_181_fu_6586_p2;
wire   [3:0] xor_ln45_138_fu_6598_p2;
wire   [3:0] xor_ln45_139_fu_6604_p2;
wire   [1:0] a1_sqr_31_fu_6639_p3;
wire   [1:0] a0_sqr_16_fu_6628_p3;
wire   [1:0] xor_ln59_16_fu_6646_p2;
wire   [1:0] a1_sqr_32_fu_6670_p3;
wire   [1:0] a0_sqr_20_fu_6663_p3;
wire   [1:0] a0_138_fu_6676_p2;
wire   [1:0] tmp_36_fu_6689_p3;
wire   [3:0] a1_sqr_33_fu_6682_p3;
wire   [3:0] a0_sqr_18_fu_6652_p3;
wire   [1:0] xor_ln28_43_fu_6695_p2;
wire   [3:0] xor_ln59_19_fu_6701_p2;
wire   [1:0] xor_ln45_183_fu_6610_p2;
wire   [7:0] tmp_37_fu_6707_p4;
wire   [7:0] tmp_35_fu_6616_p3;
wire   [5:0] tmp_113_fu_6724_p3;
wire   [5:0] tmp_112_fu_6716_p3;
wire   [5:0] xor_ln71_4_fu_6737_p2;
wire   [7:0] delta_1_fu_6731_p2;
wire   [1:0] a0_363_fu_6749_p4;
wire   [1:0] tmp_38_fu_6791_p3;
wire   [1:0] xor_ln28_45_fu_6799_p2;
wire   [1:0] a1_336_fu_6759_p4;
wire   [0:0] xor_ln70_29_fu_6819_p2;
wire   [0:0] xor_ln70_28_fu_6813_p2;
wire   [0:0] xor_ln70_32_fu_6836_p2;
wire   [0:0] xor_ln70_31_fu_6830_p2;
wire   [0:0] xor_ln70_33_fu_6842_p2;
wire   [0:0] xor_ln70_30_fu_6824_p2;
wire   [1:0] xor_ln70_36_fu_6860_p2;
wire   [1:0] xor_ln70_35_fu_6854_p2;
wire   [3:0] a0_362_fu_6743_p2;
wire   [3:0] tmp_39_fu_6805_p3;
wire   [1:0] a0_365_fu_6866_p2;
wire   [3:0] a0z1_2_fu_6872_p2;
wire   [0:0] a0_366_fu_6848_p2;
wire   [1:0] b0_53_fu_6888_p2;
wire   [0:0] a1_339_fu_6904_p3;
wire   [0:0] a_208_fu_6932_p2;
wire   [0:0] z1_53_fu_6944_p2;
wire   [0:0] z0_53_fu_6926_p2;
wire   [0:0] z2_53_fu_6950_p2;
wire   [0:0] xor_ln45_140_fu_6956_p2;
wire   [0:0] xor_ln45_141_fu_6962_p2;
wire   [1:0] a1_338_fu_6878_p4;
wire   [1:0] b1_149_fu_6894_p4;
wire   [0:0] a0_368_fu_6976_p3;
wire   [1:0] a_210_fu_6984_p2;
wire   [1:0] b_166_fu_6998_p2;
wire   [0:0] a0_367_fu_7004_p2;
wire   [0:0] a1_340_fu_7010_p3;
wire   [0:0] a_212_fu_7038_p2;
wire   [0:0] z1_54_fu_7050_p2;
wire   [0:0] z0_55_fu_7032_p2;
wire   [0:0] z2_54_fu_7056_p2;
wire   [0:0] xor_ln45_142_fu_7062_p2;
wire   [0:0] xor_ln45_143_fu_7068_p2;
wire   [0:0] a1_341_fu_7082_p3;
wire   [0:0] a_216_fu_7104_p2;
wire   [0:0] z1_56_fu_7116_p2;
wire   [0:0] z0_56_fu_7098_p2;
wire   [0:0] z2_55_fu_7122_p2;
wire   [0:0] a1_126_fu_7128_p2;
wire   [0:0] a0_150_fu_7134_p2;
wire   [0:0] xor_ln28_46_fu_7148_p2;
wire   [1:0] z1_55_fu_7074_p3;
wire   [1:0] z0_54_fu_6968_p3;
wire   [1:0] z2_191_fu_7140_p3;
wire   [1:0] tmp_40_fu_7154_p3;
wire   [1:0] xor_ln45_193_fu_7168_p2;
wire   [1:0] xor_ln45_192_fu_7162_p2;
wire   [0:0] xor_ln45_200_fu_7174_p2;
wire   [1:0] xor_ln45_148_fu_7180_p2;
wire   [1:0] xor_ln45_149_fu_7186_p2;
wire   [1:0] a1_sqr_34_fu_7236_p3;
wire   [1:0] a0_sqr_23_fu_7228_p3;
reg   [1:0] tmp_271_fu_7250_p4;
wire   [1:0] xor_ln59_21_fu_7244_p2;
wire   [0:0] xor_ln45_201_fu_7192_p2;
wire   [3:0] tmp_42_fu_7260_p3;
wire   [3:0] tmp_41_fu_7198_p3;
wire   [2:0] tmp_115_fu_7276_p3;
wire   [2:0] tmp_114_fu_7268_p3;
wire   [0:0] xor_ln36_2_fu_7302_p2;
wire   [0:0] xor_ln36_1_fu_7296_p2;
wire   [2:0] xor_ln36_fu_7290_p2;
wire   [3:0] delta_2_fu_7284_p2;
wire   [0:0] a0_372_fu_7320_p3;
wire   [0:0] a1_343_fu_7328_p3;
wire   [0:0] b_181_fu_7336_p2;
wire   [1:0] a0_371_fu_7314_p2;
wire   [1:0] tmp_43_fu_7342_p3;
wire   [0:0] a0_373_fu_7308_p2;
wire   [1:0] a0z1_3_fu_7350_p2;
wire   [0:0] b0_57_fu_7356_p2;
wire   [0:0] a1_344_fu_7362_p3;
wire   [0:0] b1_153_fu_7370_p3;
wire   [0:0] a_223_fu_7384_p2;
wire   [0:0] b_176_fu_7390_p2;
wire   [0:0] z1_57_fu_7396_p2;
wire   [0:0] z0_57_fu_7378_p2;
wire   [0:0] z2_57_fu_7402_p2;
wire   [0:0] xor_ln45_150_fu_7408_p2;
wire   [0:0] xor_ln45_151_fu_7414_p2;
wire   [1:0] tmp_45_fu_7428_p3;
wire   [1:0] tmp_44_fu_7420_p3;
wire   [1:0] delta_3_fu_7436_p2;
wire   [0:0] a0_374_fu_7442_p2;
wire   [0:0] a1_345_fu_7448_p3;
wire   [0:0] a0z1_4_fu_7456_p2;
wire   [0:0] and_ln36_fu_7462_p2;
wire   [0:0] delta_4_fu_7468_p2;
wire   [0:0] a0_375_fu_7480_p2;
wire   [0:0] a_229_fu_7492_p2;
wire   [0:0] a1_346_fu_7474_p2;
wire   [0:0] z1_58_fu_7498_p2;
wire   [0:0] z0_58_fu_7486_p2;
wire   [0:0] z2_58_fu_7504_p2;
wire   [0:0] z1_59_fu_7528_p2;
wire   [0:0] z0_59_fu_7522_p2;
wire   [0:0] z2_59_fu_7534_p2;
wire   [1:0] b_187_fu_7558_p2;
wire   [0:0] z1_60_fu_7594_p2;
wire   [0:0] z0_60_fu_7590_p2;
wire   [0:0] z2_60_fu_7598_p2;
wire   [0:0] xor_ln45_156_fu_7602_p2;
wire   [0:0] xor_ln45_157_fu_7608_p2;
wire   [1:0] a1_347_fu_7584_p3;
wire   [1:0] a0_376_fu_7578_p3;
wire   [1:0] a_235_fu_7622_p2;
wire   [0:0] a0_378_fu_7628_p2;
wire   [0:0] b0_58_fu_7640_p2;
wire   [0:0] a1_349_fu_7632_p3;
wire   [0:0] a_237_fu_7650_p2;
wire   [0:0] b_189_fu_7656_p2;
wire   [0:0] z1_61_fu_7661_p2;
wire   [0:0] z0_62_fu_7644_p2;
wire   [0:0] z2_61_fu_7667_p2;
wire   [0:0] xor_ln45_158_fu_7672_p2;
wire   [0:0] xor_ln45_159_fu_7678_p2;
wire   [0:0] z1_63_fu_7696_p2;
wire   [0:0] z0_63_fu_7692_p2;
wire   [0:0] z2_62_fu_7700_p2;
wire   [0:0] a1_141_fu_7704_p2;
wire   [0:0] a0_167_fu_7710_p2;
wire   [0:0] xor_ln28_48_fu_7724_p2;
wire   [1:0] z1_62_fu_7684_p3;
wire   [1:0] z0_61_fu_7614_p3;
wire   [1:0] z2_192_fu_7716_p3;
wire   [1:0] tmp_46_fu_7730_p3;
wire   [1:0] xor_ln45_209_fu_7744_p2;
wire   [1:0] xor_ln45_208_fu_7738_p2;
wire   [0:0] z1_64_fu_7766_p2;
wire   [0:0] z0_64_fu_7762_p2;
wire   [0:0] z2_64_fu_7770_p2;
wire   [0:0] xor_ln45_166_fu_7774_p2;
wire   [0:0] xor_ln45_167_fu_7780_p2;
wire   [0:0] z1_65_fu_7799_p2;
wire   [0:0] z0_66_fu_7794_p2;
wire   [0:0] z2_65_fu_7804_p2;
wire   [0:0] xor_ln45_168_fu_7809_p2;
wire   [0:0] xor_ln45_169_fu_7815_p2;
wire   [0:0] z1_67_fu_7833_p2;
wire   [0:0] z0_67_fu_7829_p2;
wire   [0:0] z2_66_fu_7837_p2;
wire   [0:0] a1_142_fu_7841_p2;
wire   [0:0] a0_170_fu_7847_p2;
wire   [0:0] xor_ln28_49_fu_7861_p2;
wire   [1:0] z0_65_fu_7786_p3;
wire   [1:0] z2_193_fu_7853_p3;
wire   [1:0] z1_66_fu_7821_p3;
wire   [1:0] tmp_47_fu_7867_p3;
wire   [1:0] a_250_fu_7881_p2;
wire   [1:0] a0_381_fu_7875_p2;
wire   [1:0] a1_352_fu_7887_p2;
wire   [1:0] a1_360_fu_7750_p2;
wire   [1:0] a0_389_fu_7756_p2;
wire   [0:0] a0_382_fu_7893_p2;
wire   [0:0] a1_353_fu_7915_p3;
wire   [0:0] a_248_fu_7928_p2;
wire   [0:0] z1_68_fu_7934_p2;
wire   [0:0] z0_68_fu_7923_p2;
wire   [0:0] z2_68_fu_7939_p2;
wire   [0:0] xor_ln45_176_fu_7944_p2;
wire   [0:0] xor_ln45_177_fu_7950_p2;
wire   [0:0] a0_384_fu_7964_p1;
wire   [0:0] a0_383_fu_7968_p2;
wire   [0:0] b0_60_fu_7982_p2;
wire   [0:0] a1_354_fu_7974_p3;
wire   [0:0] a_252_fu_7992_p2;
wire   [0:0] b_202_fu_7998_p2;
wire   [0:0] z1_69_fu_8003_p2;
wire   [0:0] z0_70_fu_7986_p2;
wire   [0:0] z2_69_fu_8009_p2;
wire   [0:0] xor_ln45_178_fu_8014_p2;
wire   [0:0] xor_ln45_179_fu_8020_p2;
wire   [0:0] a1_355_fu_8034_p3;
wire   [0:0] a_256_fu_8047_p2;
wire   [0:0] z1_71_fu_8053_p2;
wire   [0:0] z0_71_fu_8042_p2;
wire   [0:0] z2_70_fu_8058_p2;
wire   [0:0] a1_149_fu_8063_p2;
wire   [0:0] a0_190_fu_8069_p2;
wire   [0:0] xor_ln28_50_fu_8083_p2;
wire   [1:0] z1_70_fu_8026_p3;
wire   [1:0] z0_69_fu_7956_p3;
wire   [1:0] z2_194_fu_8075_p3;
wire   [1:0] tmp_48_fu_8089_p3;
wire   [1:0] xor_ln45_236_fu_8103_p2;
wire   [1:0] xor_ln45_235_fu_8097_p2;
wire   [1:0] xor_ln45_184_fu_8109_p2;
wire   [1:0] xor_ln45_185_fu_8115_p2;
wire   [3:0] a1_351_fu_7907_p3;
wire   [3:0] a0_380_fu_7899_p3;
wire   [3:0] a_259_fu_8133_p2;
wire   [0:0] a0_390_fu_8129_p1;
wire   [1:0] a0_385_fu_8139_p2;
wire   [0:0] a0_386_fu_8155_p2;
wire   [0:0] b0_62_fu_8169_p2;
wire   [0:0] a1_357_fu_8161_p3;
wire   [0:0] a_262_fu_8179_p2;
wire   [0:0] b_211_fu_8185_p2;
wire   [0:0] z1_72_fu_8190_p2;
wire   [0:0] z0_73_fu_8173_p2;
wire   [0:0] z2_72_fu_8196_p2;
wire   [0:0] xor_ln45_186_fu_8201_p2;
wire   [0:0] xor_ln45_187_fu_8207_p2;
wire   [1:0] a1_356_fu_8145_p4;
wire   [0:0] a0_388_fu_8221_p3;
wire   [1:0] a_264_fu_8229_p2;
wire   [0:0] a0_387_fu_8235_p2;
wire   [0:0] b0_63_fu_8249_p2;
wire   [0:0] a1_358_fu_8241_p3;
wire   [0:0] a_266_fu_8260_p2;
wire   [0:0] b_215_fu_8266_p2;
wire   [0:0] z1_73_fu_8271_p2;
wire   [0:0] z0_75_fu_8254_p2;
wire   [0:0] z2_73_fu_8277_p2;
wire   [0:0] xor_ln45_188_fu_8282_p2;
wire   [0:0] xor_ln45_189_fu_8288_p2;
wire   [0:0] a1_359_fu_8302_p3;
wire   [0:0] a_270_fu_8315_p2;
wire   [0:0] b_219_fu_8321_p2;
wire   [0:0] z1_75_fu_8325_p2;
wire   [0:0] z0_76_fu_8310_p2;
wire   [0:0] z2_74_fu_8331_p2;
wire   [0:0] a1_155_fu_8336_p2;
wire   [0:0] a0_195_fu_8342_p2;
wire   [0:0] xor_ln28_51_fu_8356_p2;
wire   [1:0] z1_74_fu_8294_p3;
wire   [1:0] z0_74_fu_8213_p3;
wire   [1:0] z2_195_fu_8348_p3;
wire   [1:0] tmp_49_fu_8362_p3;
wire   [1:0] xor_ln45_240_fu_8376_p2;
wire   [1:0] xor_ln45_239_fu_8370_p2;
wire   [1:0] xor_ln45_194_fu_8382_p2;
wire   [1:0] xor_ln45_195_fu_8388_p2;
wire   [0:0] a1_361_fu_8402_p3;
wire   [0:0] a_276_fu_8415_p2;
wire   [0:0] z1_77_fu_8421_p2;
wire   [0:0] z0_77_fu_8410_p2;
wire   [0:0] z2_76_fu_8426_p2;
wire   [0:0] xor_ln45_196_fu_8431_p2;
wire   [0:0] xor_ln45_197_fu_8437_p2;
wire   [0:0] a0_392_fu_8451_p1;
wire   [1:0] a_278_fu_8455_p2;
wire   [0:0] a0_391_fu_8461_p2;
wire   [0:0] b0_65_fu_8475_p2;
wire   [0:0] a1_362_fu_8467_p3;
wire   [0:0] a_280_fu_8485_p2;
wire   [0:0] b_228_fu_8491_p2;
wire   [0:0] z1_78_fu_8496_p2;
wire   [0:0] z0_79_fu_8479_p2;
wire   [0:0] z2_77_fu_8502_p2;
wire   [0:0] xor_ln45_198_fu_8507_p2;
wire   [0:0] xor_ln45_199_fu_8513_p2;
wire   [0:0] a1_363_fu_8527_p3;
wire   [0:0] a_284_fu_8540_p2;
wire   [0:0] z1_80_fu_8546_p2;
wire   [0:0] z0_80_fu_8535_p2;
wire   [0:0] z2_78_fu_8551_p2;
wire   [0:0] a1_161_fu_8556_p2;
wire   [0:0] a0_200_fu_8562_p2;
wire   [0:0] xor_ln28_52_fu_8576_p2;
wire   [1:0] z1_79_fu_8519_p3;
wire   [1:0] z0_78_fu_8443_p3;
wire   [1:0] z2_196_fu_8568_p3;
wire   [1:0] tmp_50_fu_8582_p3;
wire   [1:0] xor_ln45_248_fu_8596_p2;
wire   [1:0] xor_ln45_243_fu_8590_p2;
wire   [1:0] a1_364_fu_8602_p2;
wire   [1:0] a0_201_fu_8608_p2;
wire   [0:0] a0_202_fu_8622_p1;
wire   [0:0] a1_163_fu_8626_p3;
wire   [0:0] xor_ln28_53_fu_8634_p2;
wire   [1:0] tmp_51_fu_8640_p3;
wire   [1:0] xor_ln28_54_fu_8648_p2;
wire   [3:0] z1_76_fu_8394_p3;
wire   [3:0] z0_72_fu_8121_p3;
wire   [3:0] z2_197_fu_8614_p3;
wire   [3:0] tmp_52_fu_8654_p3;
wire   [3:0] xor_ln45_258_fu_8668_p2;
wire   [3:0] xor_ln45_251_fu_8662_p2;
wire   [0:0] z1_81_fu_8703_p2;
wire   [0:0] z0_81_fu_8698_p2;
wire   [0:0] z2_81_fu_8708_p2;
wire   [0:0] xor_ln45_210_fu_8713_p2;
wire   [0:0] xor_ln45_211_fu_8719_p2;
wire   [0:0] z1_82_fu_8738_p2;
wire   [0:0] z0_83_fu_8733_p2;
wire   [0:0] z2_82_fu_8743_p2;
wire   [0:0] xor_ln45_212_fu_8748_p2;
wire   [0:0] xor_ln45_213_fu_8754_p2;
wire   [0:0] z1_84_fu_8773_p2;
wire   [0:0] z0_84_fu_8768_p2;
wire   [0:0] z2_83_fu_8778_p2;
wire   [0:0] a1_164_fu_8783_p2;
wire   [0:0] a0_203_fu_8789_p2;
wire   [0:0] xor_ln28_55_fu_8803_p2;
wire   [1:0] z1_83_fu_8760_p3;
wire   [1:0] z0_82_fu_8725_p3;
wire   [1:0] z2_198_fu_8795_p3;
wire   [1:0] tmp_53_fu_8809_p3;
wire   [1:0] xor_ln45_272_fu_8823_p2;
wire   [1:0] xor_ln45_271_fu_8817_p2;
wire   [1:0] xor_ln45_218_fu_8829_p2;
wire   [1:0] xor_ln45_219_fu_8835_p2;
wire   [0:0] z1_85_fu_8854_p2;
wire   [0:0] z0_86_fu_8849_p2;
wire   [0:0] z2_85_fu_8859_p2;
wire   [0:0] xor_ln45_220_fu_8864_p2;
wire   [0:0] xor_ln45_221_fu_8870_p2;
wire   [0:0] z1_86_fu_8889_p2;
wire   [0:0] z0_88_fu_8884_p2;
wire   [0:0] z2_86_fu_8894_p2;
wire   [0:0] xor_ln45_222_fu_8899_p2;
wire   [0:0] xor_ln45_223_fu_8905_p2;
wire   [0:0] z1_88_fu_8924_p2;
wire   [0:0] z0_89_fu_8919_p2;
wire   [0:0] z2_87_fu_8929_p2;
wire   [0:0] a1_165_fu_8934_p2;
wire   [0:0] a0_204_fu_8940_p2;
wire   [0:0] xor_ln28_56_fu_8954_p2;
wire   [1:0] z1_87_fu_8911_p3;
wire   [1:0] z0_87_fu_8876_p3;
wire   [1:0] z2_199_fu_8946_p3;
wire   [1:0] tmp_54_fu_8960_p3;
wire   [1:0] xor_ln45_282_fu_8974_p2;
wire   [1:0] xor_ln45_275_fu_8968_p2;
wire   [1:0] xor_ln45_228_fu_8980_p2;
wire   [1:0] xor_ln45_229_fu_8986_p2;
wire   [0:0] z1_90_fu_9005_p2;
wire   [0:0] z0_90_fu_9000_p2;
wire   [0:0] z2_89_fu_9010_p2;
wire   [0:0] xor_ln45_230_fu_9015_p2;
wire   [0:0] xor_ln45_231_fu_9021_p2;
wire   [0:0] z1_91_fu_9040_p2;
wire   [0:0] z0_92_fu_9035_p2;
wire   [0:0] z2_90_fu_9045_p2;
wire   [0:0] xor_ln45_232_fu_9050_p2;
wire   [0:0] xor_ln45_233_fu_9056_p2;
wire   [0:0] z1_93_fu_9075_p2;
wire   [0:0] z0_93_fu_9070_p2;
wire   [0:0] z2_91_fu_9080_p2;
wire   [0:0] a1_167_fu_9085_p2;
wire   [0:0] a0_205_fu_9091_p2;
wire   [0:0] xor_ln28_57_fu_9105_p2;
wire   [1:0] z1_92_fu_9062_p3;
wire   [1:0] z0_91_fu_9027_p3;
wire   [1:0] z2_200_fu_9097_p3;
wire   [1:0] tmp_55_fu_9111_p3;
wire   [1:0] xor_ln45_292_fu_9125_p2;
wire   [1:0] xor_ln45_285_fu_9119_p2;
wire   [1:0] a1_365_fu_9131_p2;
wire   [1:0] a0_206_fu_9137_p2;
wire   [0:0] a0_207_fu_9151_p1;
wire   [0:0] a1_169_fu_9155_p3;
wire   [0:0] xor_ln28_58_fu_9163_p2;
wire   [1:0] tmp_56_fu_9169_p3;
wire   [1:0] xor_ln28_59_fu_9177_p2;
wire   [3:0] z0_85_fu_8841_p3;
wire   [3:0] z2_201_fu_9143_p3;
wire   [3:0] z1_89_fu_8992_p3;
wire   [3:0] tmp_57_fu_9183_p3;
wire   [3:0] a_309_fu_9197_p2;
wire   [3:0] a0_394_fu_9191_p2;
wire   [0:0] xor_ln43_71_fu_9227_p2;
wire   [0:0] xor_ln43_fu_9221_p2;
wire   [1:0] xor_ln45_304_fu_9209_p2;
wire   [1:0] a0_395_fu_9203_p2;
wire   [3:0] a1_367_fu_9215_p2;
wire   [1:0] xor_ln45_306_fu_9239_p2;
wire   [1:0] xor_ln45_260_fu_8680_p2;
wire   [1:0] xor_ln45_259_fu_8674_p2;
wire   [3:0] a1_395_fu_8686_p2;
wire   [3:0] a0_420_fu_8692_p2;
wire   [0:0] a0_396_fu_9233_p2;
wire   [0:0] a1_369_fu_9291_p3;
wire   [0:0] a_298_fu_9304_p2;
wire   [0:0] z1_94_fu_9310_p2;
wire   [0:0] z0_94_fu_9299_p2;
wire   [0:0] z2_94_fu_9315_p2;
wire   [0:0] xor_ln45_244_fu_9320_p2;
wire   [0:0] xor_ln45_245_fu_9326_p2;
wire   [1:0] a1_368_fu_9281_p4;
wire   [0:0] a0_398_fu_9340_p3;
wire   [1:0] a_300_fu_9348_p2;
wire   [0:0] a0_397_fu_9354_p2;
wire   [0:0] b0_68_fu_9368_p2;
wire   [0:0] a1_370_fu_9360_p3;
wire   [0:0] a_302_fu_9378_p2;
wire   [0:0] b_242_fu_9384_p2;
wire   [0:0] z1_95_fu_9389_p2;
wire   [0:0] z0_96_fu_9372_p2;
wire   [0:0] z2_95_fu_9395_p2;
wire   [0:0] xor_ln45_246_fu_9400_p2;
wire   [0:0] xor_ln45_247_fu_9406_p2;
wire   [0:0] a1_371_fu_9420_p3;
wire   [0:0] a_306_fu_9433_p2;
wire   [0:0] z1_97_fu_9439_p2;
wire   [0:0] z0_97_fu_9428_p2;
wire   [0:0] z2_96_fu_9444_p2;
wire   [0:0] a1_178_fu_9449_p2;
wire   [0:0] a0_214_fu_9455_p2;
wire   [0:0] xor_ln28_60_fu_9469_p2;
wire   [1:0] z1_96_fu_9412_p3;
wire   [1:0] z0_95_fu_9332_p3;
wire   [1:0] z2_202_fu_9461_p3;
wire   [1:0] tmp_58_fu_9475_p3;
wire   [1:0] xor_ln45_316_fu_9489_p2;
wire   [1:0] xor_ln45_309_fu_9483_p2;
wire   [1:0] xor_ln45_252_fu_9495_p2;
wire   [1:0] xor_ln45_253_fu_9501_p2;
wire   [1:0] a0_403_fu_9519_p1;
wire   [0:0] a0_404_fu_9515_p1;
wire   [1:0] a0_399_fu_9523_p2;
wire   [0:0] a0_400_fu_9539_p2;
wire   [0:0] b0_70_fu_9553_p2;
wire   [0:0] a1_373_fu_9545_p3;
wire   [0:0] a_312_fu_9563_p2;
wire   [0:0] b_251_fu_9569_p2;
wire   [0:0] z1_98_fu_9574_p2;
wire   [0:0] z0_99_fu_9557_p2;
wire   [0:0] z2_98_fu_9580_p2;
wire   [0:0] xor_ln45_254_fu_9585_p2;
wire   [0:0] xor_ln45_255_fu_9591_p2;
wire   [1:0] a1_372_fu_9529_p4;
wire   [0:0] a0_402_fu_9605_p3;
wire   [1:0] a_314_fu_9613_p2;
wire   [0:0] a0_401_fu_9619_p2;
wire   [0:0] b0_71_fu_9633_p2;
wire   [0:0] a1_374_fu_9625_p3;
wire   [0:0] a_316_fu_9644_p2;
wire   [0:0] b_255_fu_9650_p2;
wire   [0:0] z1_99_fu_9655_p2;
wire   [0:0] z0_101_fu_9638_p2;
wire   [0:0] z2_99_fu_9661_p2;
wire   [0:0] xor_ln45_256_fu_9666_p2;
wire   [0:0] xor_ln45_257_fu_9672_p2;
wire   [0:0] a1_375_fu_9686_p3;
wire   [0:0] a_320_fu_9699_p2;
wire   [0:0] b_259_fu_9705_p2;
wire   [0:0] z1_101_fu_9709_p2;
wire   [0:0] z0_102_fu_9694_p2;
wire   [0:0] z2_100_fu_9715_p2;
wire   [0:0] a1_183_fu_9720_p2;
wire   [0:0] a0_219_fu_9726_p2;
wire   [0:0] xor_ln28_61_fu_9740_p2;
wire   [1:0] z1_100_fu_9678_p3;
wire   [1:0] z0_100_fu_9597_p3;
wire   [1:0] z2_203_fu_9732_p3;
wire   [1:0] tmp_59_fu_9746_p3;
wire   [1:0] xor_ln45_326_fu_9760_p2;
wire   [1:0] xor_ln45_319_fu_9754_p2;
wire   [1:0] xor_ln45_262_fu_9766_p2;
wire   [1:0] xor_ln45_263_fu_9772_p2;
wire   [0:0] a1_377_fu_9796_p3;
wire   [0:0] a_326_fu_9809_p2;
wire   [0:0] z1_103_fu_9815_p2;
wire   [0:0] z0_103_fu_9804_p2;
wire   [0:0] z2_102_fu_9820_p2;
wire   [0:0] xor_ln45_264_fu_9825_p2;
wire   [0:0] xor_ln45_265_fu_9831_p2;
wire   [1:0] a1_376_fu_9786_p4;
wire   [0:0] a0_406_fu_9845_p3;
wire   [1:0] a_328_fu_9853_p2;
wire   [0:0] a0_405_fu_9859_p2;
wire   [0:0] b0_74_fu_9873_p2;
wire   [0:0] a1_378_fu_9865_p3;
wire   [0:0] a_330_fu_9883_p2;
wire   [0:0] b_268_fu_9889_p2;
wire   [0:0] z1_104_fu_9894_p2;
wire   [0:0] z0_105_fu_9877_p2;
wire   [0:0] z2_103_fu_9900_p2;
wire   [0:0] xor_ln45_266_fu_9905_p2;
wire   [0:0] xor_ln45_267_fu_9911_p2;
wire   [0:0] a1_379_fu_9925_p3;
wire   [0:0] a_334_fu_9938_p2;
wire   [0:0] z1_106_fu_9944_p2;
wire   [0:0] z0_106_fu_9933_p2;
wire   [0:0] z2_104_fu_9949_p2;
wire   [0:0] a1_190_fu_9954_p2;
wire   [0:0] a0_224_fu_9960_p2;
wire   [0:0] xor_ln28_62_fu_9974_p2;
wire   [1:0] z1_105_fu_9917_p3;
wire   [1:0] z0_104_fu_9837_p3;
wire   [1:0] z2_204_fu_9966_p3;
wire   [1:0] tmp_60_fu_9980_p3;
wire   [1:0] xor_ln45_336_fu_9994_p2;
wire   [1:0] xor_ln45_329_fu_9988_p2;
wire   [1:0] a1_380_fu_10000_p2;
wire   [1:0] a0_225_fu_10006_p2;
wire   [0:0] a0_226_fu_10020_p1;
wire   [0:0] a1_192_fu_10024_p3;
wire   [0:0] xor_ln28_63_fu_10032_p2;
wire   [1:0] tmp_61_fu_10038_p3;
wire   [1:0] xor_ln28_64_fu_10046_p2;
wire   [3:0] z1_102_fu_9778_p3;
wire   [3:0] z0_98_fu_9507_p3;
wire   [3:0] z2_205_fu_10012_p3;
wire   [3:0] tmp_62_fu_10052_p3;
wire   [3:0] xor_ln45_340_fu_10066_p2;
wire   [3:0] xor_ln45_339_fu_10060_p2;
wire   [3:0] xor_ln45_276_fu_10072_p2;
wire   [3:0] xor_ln45_277_fu_10078_p2;
wire   [1:0] a0_429_fu_10100_p1;
wire   [7:0] a1_366_fu_9273_p3;
wire   [7:0] a0_393_fu_9245_p3;
wire   [5:0] trunc_ln43_2_fu_10104_p3;
wire   [5:0] a0_419_cast_fu_9253_p3;
wire   [7:0] a_339_fu_10112_p2;
wire   [1:0] a0_421_fu_10096_p1;
wire   [3:0] a0_407_fu_10124_p2;
wire   [0:0] a0_422_fu_10092_p1;
wire   [1:0] a0_408_fu_10140_p2;
wire   [0:0] a0_409_fu_10156_p2;
wire   [0:0] b0_77_fu_10170_p2;
wire   [0:0] a1_383_fu_10162_p3;
wire   [0:0] a_343_fu_10180_p2;
wire   [0:0] b_278_fu_10186_p2;
wire   [0:0] z1_107_fu_10191_p2;
wire   [0:0] z0_108_fu_10174_p2;
wire   [0:0] z2_107_fu_10197_p2;
wire   [0:0] xor_ln45_278_fu_10202_p2;
wire   [0:0] xor_ln45_279_fu_10208_p2;
wire   [1:0] a1_382_fu_10146_p4;
wire   [0:0] a0_411_fu_10222_p3;
wire   [1:0] a_345_fu_10230_p2;
wire   [0:0] a0_410_fu_10236_p2;
wire   [0:0] b0_78_fu_10250_p2;
wire   [0:0] a1_384_fu_10242_p3;
wire   [0:0] a_347_fu_10261_p2;
wire   [0:0] b_282_fu_10267_p2;
wire   [0:0] z1_108_fu_10272_p2;
wire   [0:0] z0_110_fu_10255_p2;
wire   [0:0] z2_108_fu_10278_p2;
wire   [0:0] xor_ln45_280_fu_10283_p2;
wire   [0:0] xor_ln45_281_fu_10289_p2;
wire   [0:0] a1_385_fu_10303_p3;
wire   [0:0] a_351_fu_10316_p2;
wire   [0:0] b_286_fu_10322_p2;
wire   [0:0] z1_110_fu_10326_p2;
wire   [0:0] z0_111_fu_10311_p2;
wire   [0:0] z2_109_fu_10332_p2;
wire   [0:0] a1_198_fu_10337_p2;
wire   [0:0] a0_232_fu_10343_p2;
wire   [0:0] xor_ln28_65_fu_10357_p2;
wire   [1:0] z1_109_fu_10295_p3;
wire   [1:0] z0_109_fu_10214_p3;
wire   [1:0] z2_206_fu_10349_p3;
wire   [1:0] tmp_63_fu_10363_p3;
wire   [1:0] xor_ln45_344_fu_10377_p2;
wire   [1:0] xor_ln45_343_fu_10371_p2;
wire   [1:0] xor_ln45_286_fu_10383_p2;
wire   [1:0] xor_ln45_287_fu_10389_p2;
wire   [3:0] a1_381_fu_10130_p4;
wire   [1:0] a0_416_fu_10411_p4;
wire   [3:0] a_354_fu_10421_p2;
wire   [0:0] a0_417_fu_10403_p3;
wire   [1:0] a0_412_fu_10427_p2;
wire   [0:0] a0_413_fu_10443_p2;
wire   [0:0] b0_81_fu_10457_p2;
wire   [0:0] a1_387_fu_10449_p3;
wire   [0:0] a_357_fu_10468_p2;
wire   [0:0] b_291_fu_10474_p2;
wire   [0:0] z1_111_fu_10479_p2;
wire   [0:0] z0_113_fu_10462_p2;
wire   [0:0] z2_111_fu_10485_p2;
wire   [0:0] xor_ln45_288_fu_10490_p2;
wire   [0:0] xor_ln45_289_fu_10496_p2;
wire   [1:0] a1_386_fu_10433_p4;
wire   [0:0] a0_415_fu_10510_p3;
wire   [1:0] a_359_fu_10518_p2;
wire   [0:0] a0_414_fu_10524_p2;
wire   [0:0] b0_82_fu_10538_p2;
wire   [0:0] a1_388_fu_10530_p3;
wire   [0:0] a_361_fu_10549_p2;
wire   [0:0] b_295_fu_10555_p2;
wire   [0:0] z1_112_fu_10560_p2;
wire   [0:0] z0_115_fu_10543_p2;
wire   [0:0] z2_112_fu_10566_p2;
wire   [0:0] xor_ln45_290_fu_10571_p2;
wire   [0:0] xor_ln45_291_fu_10577_p2;
wire   [0:0] a1_389_fu_10591_p3;
wire   [0:0] a_365_fu_10604_p2;
wire   [0:0] b_299_fu_10610_p2;
wire   [0:0] z1_114_fu_10614_p2;
wire   [0:0] z0_116_fu_10599_p2;
wire   [0:0] z2_113_fu_10620_p2;
wire   [0:0] a1_212_fu_10625_p2;
wire   [0:0] a0_237_fu_10631_p2;
wire   [0:0] xor_ln28_66_fu_10645_p2;
wire   [1:0] z1_113_fu_10583_p3;
wire   [1:0] z0_114_fu_10502_p3;
wire   [1:0] z2_207_fu_10637_p3;
wire   [1:0] tmp_64_fu_10651_p3;
wire   [1:0] xor_ln45_354_fu_10665_p2;
wire   [1:0] xor_ln45_347_fu_10659_p2;
wire   [1:0] xor_ln45_296_fu_10671_p2;
wire   [1:0] xor_ln45_297_fu_10677_p2;
wire   [5:0] xor_ln43_83_fu_10118_p2;
wire   [0:0] a1_391_fu_10701_p3;
wire   [0:0] a_371_fu_10714_p2;
wire   [0:0] b_304_fu_10720_p2;
wire   [0:0] z1_116_fu_10724_p2;
wire   [0:0] z0_117_fu_10709_p2;
wire   [0:0] z2_115_fu_10730_p2;
wire   [0:0] xor_ln45_298_fu_10735_p2;
wire   [0:0] xor_ln45_299_fu_10741_p2;
wire   [1:0] a1_390_fu_10691_p4;
wire   [0:0] a0_419_fu_10755_p3;
wire   [1:0] a_373_fu_10763_p2;
wire   [0:0] a0_418_fu_10769_p2;
wire   [0:0] b0_86_fu_10783_p2;
wire   [0:0] a1_392_fu_10775_p3;
wire   [0:0] a_375_fu_10793_p2;
wire   [0:0] b_308_fu_10799_p2;
wire   [0:0] z1_117_fu_10804_p2;
wire   [0:0] z0_119_fu_10787_p2;
wire   [0:0] z2_116_fu_10810_p2;
wire   [0:0] xor_ln45_300_fu_10815_p2;
wire   [0:0] xor_ln45_301_fu_10821_p2;
wire   [0:0] a1_393_fu_10835_p3;
wire   [0:0] a_379_fu_10848_p2;
wire   [0:0] b_312_fu_10854_p2;
wire   [0:0] z1_119_fu_10858_p2;
wire   [0:0] z0_120_fu_10843_p2;
wire   [0:0] z2_117_fu_10864_p2;
wire   [0:0] a1_217_fu_10869_p2;
wire   [0:0] a0_242_fu_10875_p2;
wire   [0:0] xor_ln28_67_fu_10889_p2;
wire   [1:0] z1_118_fu_10827_p3;
wire   [1:0] z0_118_fu_10747_p3;
wire   [1:0] z2_208_fu_10881_p3;
wire   [1:0] tmp_65_fu_10895_p3;
wire   [1:0] xor_ln45_364_fu_10909_p2;
wire   [1:0] xor_ln45_357_fu_10903_p2;
wire   [1:0] a1_394_fu_10915_p2;
wire   [1:0] a0_243_fu_10921_p2;
wire   [0:0] a0_244_fu_10935_p1;
wire   [0:0] a1_219_fu_10939_p3;
wire   [0:0] xor_ln28_68_fu_10947_p2;
wire   [1:0] tmp_66_fu_10953_p3;
wire   [1:0] xor_ln28_69_fu_10961_p2;
wire   [3:0] z1_115_fu_10683_p3;
wire   [3:0] z0_112_fu_10395_p3;
wire   [3:0] z2_209_fu_10927_p3;
wire   [3:0] tmp_67_fu_10967_p3;
wire   [3:0] xor_ln45_374_fu_10981_p2;
wire   [3:0] xor_ln45_367_fu_10975_p2;
wire   [3:0] xor_ln45_310_fu_10987_p2;
wire   [3:0] xor_ln45_311_fu_10993_p2;
wire   [1:0] xor_ln73_fu_9261_p2;
wire   [0:0] a1_397_fu_11017_p3;
wire   [0:0] a_388_fu_11030_p2;
wire   [0:0] z1_121_fu_11036_p2;
wire   [0:0] z0_121_fu_11025_p2;
wire   [0:0] z2_120_fu_11041_p2;
wire   [0:0] xor_ln45_312_fu_11046_p2;
wire   [0:0] xor_ln45_313_fu_11052_p2;
wire   [1:0] a1_396_fu_11007_p4;
wire   [0:0] a0_424_fu_11066_p3;
wire   [1:0] a_390_fu_11074_p2;
wire   [0:0] a0_423_fu_11080_p2;
wire   [0:0] b0_89_fu_11094_p2;
wire   [0:0] a1_398_fu_11086_p3;
wire   [0:0] a_392_fu_11104_p2;
wire   [0:0] b_322_fu_11110_p2;
wire   [0:0] z1_122_fu_11115_p2;
wire   [0:0] z0_123_fu_11098_p2;
wire   [0:0] z2_121_fu_11121_p2;
wire   [0:0] xor_ln45_314_fu_11126_p2;
wire   [0:0] xor_ln45_315_fu_11132_p2;
wire   [0:0] a1_399_fu_11146_p3;
wire   [0:0] a_396_fu_11159_p2;
wire   [0:0] z1_124_fu_11165_p2;
wire   [0:0] z0_124_fu_11154_p2;
wire   [0:0] z2_122_fu_11170_p2;
wire   [0:0] a1_225_fu_11175_p2;
wire   [0:0] a0_250_fu_11181_p2;
wire   [0:0] xor_ln28_70_fu_11195_p2;
wire   [1:0] z1_123_fu_11138_p3;
wire   [1:0] z0_122_fu_11058_p3;
wire   [1:0] z2_210_fu_11187_p3;
wire   [1:0] tmp_68_fu_11201_p3;
wire   [1:0] xor_ln45_378_fu_11215_p2;
wire   [1:0] xor_ln45_377_fu_11209_p2;
wire   [1:0] xor_ln45_320_fu_11221_p2;
wire   [1:0] xor_ln45_321_fu_11227_p2;
wire   [3:0] a_399_fu_11245_p2;
wire   [0:0] a0_430_fu_11241_p1;
wire   [1:0] a0_425_fu_11251_p2;
wire   [0:0] a0_426_fu_11267_p2;
wire   [0:0] b0_91_fu_11281_p2;
wire   [0:0] a1_401_fu_11273_p3;
wire   [0:0] a_402_fu_11291_p2;
wire   [0:0] b_331_fu_11297_p2;
wire   [0:0] z1_125_fu_11302_p2;
wire   [0:0] z0_126_fu_11285_p2;
wire   [0:0] z2_124_fu_11308_p2;
wire   [0:0] xor_ln45_322_fu_11313_p2;
wire   [0:0] xor_ln45_323_fu_11319_p2;
wire   [1:0] a1_400_fu_11257_p4;
wire   [0:0] a0_428_fu_11333_p3;
wire   [1:0] a_404_fu_11341_p2;
wire   [0:0] a0_427_fu_11347_p2;
wire   [0:0] b0_92_fu_11361_p2;
wire   [0:0] a1_402_fu_11353_p3;
wire   [0:0] a_406_fu_11372_p2;
wire   [0:0] b_335_fu_11378_p2;
wire   [0:0] z1_126_fu_11383_p2;
wire   [0:0] z0_128_fu_11366_p2;
wire   [0:0] z2_125_fu_11389_p2;
wire   [0:0] xor_ln45_324_fu_11394_p2;
wire   [0:0] xor_ln45_325_fu_11400_p2;
wire   [0:0] a1_403_fu_11414_p3;
wire   [0:0] a_410_fu_11427_p2;
wire   [0:0] b_339_fu_11433_p2;
wire   [0:0] z1_128_fu_11437_p2;
wire   [0:0] z0_129_fu_11422_p2;
wire   [0:0] z2_126_fu_11443_p2;
wire   [0:0] a1_230_fu_11448_p2;
wire   [0:0] a0_255_fu_11454_p2;
wire   [0:0] xor_ln28_71_fu_11468_p2;
wire   [1:0] z1_127_fu_11406_p3;
wire   [1:0] z0_127_fu_11325_p3;
wire   [1:0] z2_211_fu_11460_p3;
wire   [1:0] tmp_69_fu_11474_p3;
wire   [1:0] xor_ln45_388_fu_11488_p2;
wire   [1:0] xor_ln45_381_fu_11482_p2;
wire   [1:0] xor_ln45_330_fu_11494_p2;
wire   [1:0] xor_ln45_331_fu_11500_p2;
wire   [1:0] xor_ln73_1_fu_9267_p2;
wire   [0:0] a1_405_fu_11524_p3;
wire   [0:0] a_416_fu_11537_p2;
wire   [0:0] z1_130_fu_11543_p2;
wire   [0:0] z0_130_fu_11532_p2;
wire   [0:0] z2_128_fu_11548_p2;
wire   [0:0] xor_ln45_332_fu_11553_p2;
wire   [0:0] xor_ln45_333_fu_11559_p2;
wire   [1:0] a1_404_fu_11514_p4;
wire   [0:0] a0_432_fu_11573_p3;
wire   [1:0] a_418_fu_11581_p2;
wire   [0:0] a0_431_fu_11587_p2;
wire   [0:0] b0_94_fu_11601_p2;
wire   [0:0] a1_406_fu_11593_p3;
wire   [0:0] a_420_fu_11611_p2;
wire   [0:0] b_348_fu_11617_p2;
wire   [0:0] z1_131_fu_11622_p2;
wire   [0:0] z0_132_fu_11605_p2;
wire   [0:0] z2_129_fu_11628_p2;
wire   [0:0] xor_ln45_334_fu_11633_p2;
wire   [0:0] xor_ln45_335_fu_11639_p2;
wire   [0:0] a1_407_fu_11653_p3;
wire   [0:0] a_424_fu_11666_p2;
wire   [0:0] z1_133_fu_11672_p2;
wire   [0:0] z0_133_fu_11661_p2;
wire   [0:0] z2_130_fu_11677_p2;
wire   [0:0] a1_fu_11682_p2;
wire   [0:0] a0_260_fu_11688_p2;
wire   [0:0] xor_ln28_fu_11702_p2;
wire   [1:0] z1_132_fu_11645_p3;
wire   [1:0] z0_131_fu_11565_p3;
wire   [1:0] z2_212_fu_11694_p3;
wire   [1:0] tmp_70_fu_11708_p3;
wire   [1:0] xor_ln45_398_fu_11722_p2;
wire   [1:0] xor_ln45_391_fu_11716_p2;
wire   [1:0] a1_408_fu_11728_p2;
wire   [1:0] a0_261_fu_11734_p2;
wire   [0:0] a0_262_fu_11748_p1;
wire   [0:0] a1_236_fu_11752_p3;
wire   [0:0] xor_ln28_72_fu_11760_p2;
wire   [1:0] tmp_71_fu_11766_p3;
wire   [1:0] xor_ln28_73_fu_11774_p2;
wire   [3:0] z1_129_fu_11506_p3;
wire   [3:0] z0_125_fu_11233_p3;
wire   [3:0] z2_213_fu_11740_p3;
wire   [3:0] tmp_72_fu_11780_p3;
wire   [3:0] xor_ln45_408_fu_11794_p2;
wire   [3:0] xor_ln45_401_fu_11788_p2;
wire   [3:0] a1_409_fu_11800_p2;
wire   [3:0] a0_263_fu_11806_p2;
wire   [0:0] a0_265_fu_11834_p3;
wire   [0:0] a1_239_fu_11842_p3;
wire   [0:0] xor_ln28_74_fu_11850_p2;
wire   [1:0] a0_264_fu_11820_p1;
wire   [1:0] tmp_73_fu_11856_p3;
wire   [1:0] xor_ln28_75_fu_11864_p2;
wire   [1:0] a1_410_fu_11824_p4;
wire   [3:0] tmp_74_fu_11870_p3;
wire   [3:0] xor_ln28_76_fu_11878_p2;
wire   [7:0] z1_120_fu_10999_p3;
wire   [7:0] z0_107_fu_10084_p3;
wire   [7:0] z2_214_fu_11812_p3;
wire   [7:0] tmp_75_fu_11884_p3;
wire   [7:0] xor_ln45_412_fu_11898_p2;
wire   [7:0] xor_ln45_411_fu_11892_p2;
wire   [0:0] z1_134_fu_11921_p2;
wire   [0:0] z0_134_fu_11916_p2;
wire   [0:0] z2_134_fu_11926_p2;
wire   [0:0] xor_ln45_350_fu_11931_p2;
wire   [0:0] xor_ln45_351_fu_11937_p2;
wire   [0:0] z1_135_fu_11956_p2;
wire   [0:0] z0_136_fu_11951_p2;
wire   [0:0] z2_135_fu_11961_p2;
wire   [0:0] xor_ln45_352_fu_11966_p2;
wire   [0:0] xor_ln45_353_fu_11972_p2;
wire   [0:0] z1_137_fu_11991_p2;
wire   [0:0] z0_137_fu_11986_p2;
wire   [0:0] z2_136_fu_11996_p2;
wire   [0:0] a1_240_fu_12001_p2;
wire   [0:0] a0_266_fu_12007_p2;
wire   [0:0] xor_ln28_77_fu_12021_p2;
wire   [1:0] z1_136_fu_11978_p3;
wire   [1:0] z0_135_fu_11943_p3;
wire   [1:0] z2_215_fu_12013_p3;
wire   [1:0] tmp_76_fu_12027_p3;
wire   [1:0] xor_ln45_422_fu_12041_p2;
wire   [1:0] xor_ln45_415_fu_12035_p2;
wire   [1:0] xor_ln45_358_fu_12047_p2;
wire   [1:0] xor_ln45_359_fu_12053_p2;
wire   [0:0] z1_138_fu_12072_p2;
wire   [0:0] z0_139_fu_12067_p2;
wire   [0:0] z2_138_fu_12077_p2;
wire   [0:0] xor_ln45_360_fu_12082_p2;
wire   [0:0] xor_ln45_361_fu_12088_p2;
wire   [0:0] z1_139_fu_12107_p2;
wire   [0:0] z0_141_fu_12102_p2;
wire   [0:0] z2_139_fu_12112_p2;
wire   [0:0] xor_ln45_362_fu_12117_p2;
wire   [0:0] xor_ln45_363_fu_12123_p2;
wire   [0:0] z1_141_fu_12142_p2;
wire   [0:0] z0_142_fu_12137_p2;
wire   [0:0] z2_140_fu_12147_p2;
wire   [0:0] a1_241_fu_12152_p2;
wire   [0:0] a0_267_fu_12158_p2;
wire   [0:0] xor_ln28_78_fu_12172_p2;
wire   [1:0] z1_140_fu_12129_p3;
wire   [1:0] z0_140_fu_12094_p3;
wire   [1:0] z2_216_fu_12164_p3;
wire   [1:0] tmp_77_fu_12178_p3;
wire   [1:0] xor_ln45_432_fu_12192_p2;
wire   [1:0] xor_ln45_425_fu_12186_p2;
wire   [1:0] xor_ln45_368_fu_12198_p2;
wire   [1:0] xor_ln45_369_fu_12204_p2;
wire   [0:0] z1_143_fu_12223_p2;
wire   [0:0] z0_143_fu_12218_p2;
wire   [0:0] z2_142_fu_12228_p2;
wire   [0:0] xor_ln45_370_fu_12233_p2;
wire   [0:0] xor_ln45_371_fu_12239_p2;
wire   [0:0] z1_144_fu_12258_p2;
wire   [0:0] z0_145_fu_12253_p2;
wire   [0:0] z2_143_fu_12263_p2;
wire   [0:0] xor_ln45_372_fu_12268_p2;
wire   [0:0] xor_ln45_373_fu_12274_p2;
wire   [0:0] z1_146_fu_12293_p2;
wire   [0:0] z0_146_fu_12288_p2;
wire   [0:0] z2_144_fu_12298_p2;
wire   [0:0] a1_242_fu_12303_p2;
wire   [0:0] a0_268_fu_12309_p2;
wire   [0:0] xor_ln28_79_fu_12323_p2;
wire   [1:0] z1_145_fu_12280_p3;
wire   [1:0] z0_144_fu_12245_p3;
wire   [1:0] z2_217_fu_12315_p3;
wire   [1:0] tmp_78_fu_12329_p3;
wire   [1:0] xor_ln45_442_fu_12343_p2;
wire   [1:0] xor_ln45_435_fu_12337_p2;
wire   [1:0] a1_411_fu_12349_p2;
wire   [1:0] a0_269_fu_12355_p2;
wire   [0:0] a0_270_fu_12369_p1;
wire   [0:0] a1_244_fu_12373_p3;
wire   [0:0] xor_ln28_80_fu_12381_p2;
wire   [1:0] tmp_79_fu_12387_p3;
wire   [1:0] xor_ln28_81_fu_12395_p2;
wire   [3:0] z1_142_fu_12210_p3;
wire   [3:0] z0_138_fu_12059_p3;
wire   [3:0] z2_218_fu_12361_p3;
wire   [3:0] tmp_80_fu_12401_p3;
wire   [3:0] xor_ln45_446_fu_12415_p2;
wire   [3:0] xor_ln45_445_fu_12409_p2;
wire   [3:0] xor_ln45_382_fu_12421_p2;
wire   [3:0] xor_ln45_383_fu_12427_p2;
wire   [0:0] z1_147_fu_12446_p2;
wire   [0:0] z0_148_fu_12441_p2;
wire   [0:0] z2_147_fu_12451_p2;
wire   [0:0] xor_ln45_384_fu_12456_p2;
wire   [0:0] xor_ln45_385_fu_12462_p2;
wire   [0:0] z1_148_fu_12481_p2;
wire   [0:0] z0_150_fu_12476_p2;
wire   [0:0] z2_148_fu_12486_p2;
wire   [0:0] xor_ln45_386_fu_12491_p2;
wire   [0:0] xor_ln45_387_fu_12497_p2;
wire   [0:0] z1_150_fu_12516_p2;
wire   [0:0] z0_151_fu_12511_p2;
wire   [0:0] z2_149_fu_12521_p2;
wire   [0:0] a1_245_fu_12526_p2;
wire   [0:0] a0_271_fu_12532_p2;
wire   [0:0] xor_ln28_82_fu_12546_p2;
wire   [1:0] z1_149_fu_12503_p3;
wire   [1:0] z0_149_fu_12468_p3;
wire   [1:0] z2_219_fu_12538_p3;
wire   [1:0] tmp_81_fu_12552_p3;
wire   [1:0] xor_ln45_450_fu_12566_p2;
wire   [1:0] xor_ln45_449_fu_12560_p2;
wire   [1:0] xor_ln45_392_fu_12572_p2;
wire   [1:0] xor_ln45_393_fu_12578_p2;
wire   [0:0] z1_151_fu_12597_p2;
wire   [0:0] z0_153_fu_12592_p2;
wire   [0:0] z2_151_fu_12602_p2;
wire   [0:0] xor_ln45_394_fu_12607_p2;
wire   [0:0] xor_ln45_395_fu_12613_p2;
wire   [0:0] z1_152_fu_12632_p2;
wire   [0:0] z0_155_fu_12627_p2;
wire   [0:0] z2_152_fu_12637_p2;
wire   [0:0] xor_ln45_396_fu_12642_p2;
wire   [0:0] xor_ln45_397_fu_12648_p2;
wire   [0:0] z1_154_fu_12667_p2;
wire   [0:0] z0_156_fu_12662_p2;
wire   [0:0] z2_153_fu_12672_p2;
wire   [0:0] a1_246_fu_12677_p2;
wire   [0:0] a0_272_fu_12683_p2;
wire   [0:0] xor_ln28_83_fu_12697_p2;
wire   [1:0] z1_153_fu_12654_p3;
wire   [1:0] z0_154_fu_12619_p3;
wire   [1:0] z2_220_fu_12689_p3;
wire   [1:0] tmp_82_fu_12703_p3;
wire   [1:0] xor_ln45_456_fu_12717_p2;
wire   [1:0] xor_ln45_453_fu_12711_p2;
wire   [1:0] xor_ln45_402_fu_12723_p2;
wire   [1:0] xor_ln45_403_fu_12729_p2;
wire   [0:0] z1_156_fu_12748_p2;
wire   [0:0] z0_157_fu_12743_p2;
wire   [0:0] z2_155_fu_12753_p2;
wire   [0:0] xor_ln45_404_fu_12758_p2;
wire   [0:0] xor_ln45_405_fu_12764_p2;
wire   [0:0] z1_157_fu_12783_p2;
wire   [0:0] z0_159_fu_12778_p2;
wire   [0:0] z2_156_fu_12788_p2;
wire   [0:0] xor_ln45_406_fu_12793_p2;
wire   [0:0] xor_ln45_407_fu_12799_p2;
wire   [0:0] z1_159_fu_12818_p2;
wire   [0:0] z0_160_fu_12813_p2;
wire   [0:0] z2_157_fu_12823_p2;
wire   [0:0] a1_247_fu_12828_p2;
wire   [0:0] a0_273_fu_12834_p2;
wire   [0:0] xor_ln28_84_fu_12848_p2;
wire   [1:0] z1_158_fu_12805_p3;
wire   [1:0] z0_158_fu_12770_p3;
wire   [1:0] z2_221_fu_12840_p3;
wire   [1:0] tmp_83_fu_12854_p3;
wire   [1:0] xor_ln45_460_fu_12868_p2;
wire   [1:0] xor_ln45_459_fu_12862_p2;
wire   [1:0] a1_412_fu_12874_p2;
wire   [1:0] a0_274_fu_12880_p2;
wire   [0:0] a0_275_fu_12894_p1;
wire   [0:0] a1_249_fu_12898_p3;
wire   [0:0] xor_ln28_85_fu_12906_p2;
wire   [1:0] tmp_84_fu_12912_p3;
wire   [1:0] xor_ln28_86_fu_12920_p2;
wire   [3:0] z1_155_fu_12735_p3;
wire   [3:0] z0_152_fu_12584_p3;
wire   [3:0] z2_222_fu_12886_p3;
wire   [3:0] tmp_85_fu_12926_p3;
wire   [3:0] xor_ln45_464_fu_12940_p2;
wire   [3:0] xor_ln45_463_fu_12934_p2;
wire   [3:0] xor_ln45_416_fu_12946_p2;
wire   [3:0] xor_ln45_417_fu_12952_p2;
wire   [0:0] z1_161_fu_12971_p2;
wire   [0:0] z0_161_fu_12966_p2;
wire   [0:0] z2_160_fu_12976_p2;
wire   [0:0] xor_ln45_418_fu_12981_p2;
wire   [0:0] xor_ln45_419_fu_12987_p2;
wire   [0:0] z1_162_fu_13006_p2;
wire   [0:0] z0_163_fu_13001_p2;
wire   [0:0] z2_161_fu_13011_p2;
wire   [0:0] xor_ln45_420_fu_13016_p2;
wire   [0:0] xor_ln45_421_fu_13022_p2;
wire   [0:0] z1_164_fu_13041_p2;
wire   [0:0] z0_164_fu_13036_p2;
wire   [0:0] z2_162_fu_13046_p2;
wire   [0:0] a1_250_fu_13051_p2;
wire   [0:0] a0_276_fu_13057_p2;
wire   [0:0] xor_ln28_87_fu_13071_p2;
wire   [1:0] z1_163_fu_13028_p3;
wire   [1:0] z0_162_fu_12993_p3;
wire   [1:0] z2_223_fu_13063_p3;
wire   [1:0] tmp_86_fu_13077_p3;
wire   [1:0] xor_ln45_468_fu_13091_p2;
wire   [1:0] xor_ln45_467_fu_13085_p2;
wire   [1:0] xor_ln45_426_fu_13097_p2;
wire   [1:0] xor_ln45_427_fu_13103_p2;
wire   [0:0] z1_165_fu_13122_p2;
wire   [0:0] z0_166_fu_13117_p2;
wire   [0:0] z2_164_fu_13127_p2;
wire   [0:0] xor_ln45_428_fu_13132_p2;
wire   [0:0] xor_ln45_429_fu_13138_p2;
wire   [0:0] z1_166_fu_13157_p2;
wire   [0:0] z0_168_fu_13152_p2;
wire   [0:0] z2_165_fu_13162_p2;
wire   [0:0] xor_ln45_430_fu_13167_p2;
wire   [0:0] xor_ln45_431_fu_13173_p2;
wire   [0:0] z1_168_fu_13192_p2;
wire   [0:0] z0_169_fu_13187_p2;
wire   [0:0] z2_166_fu_13197_p2;
wire   [0:0] a1_251_fu_13202_p2;
wire   [0:0] a0_277_fu_13208_p2;
wire   [0:0] xor_ln28_88_fu_13222_p2;
wire   [1:0] z1_167_fu_13179_p3;
wire   [1:0] z0_167_fu_13144_p3;
wire   [1:0] z2_224_fu_13214_p3;
wire   [1:0] tmp_87_fu_13228_p3;
wire   [1:0] xor_ln45_472_fu_13242_p2;
wire   [1:0] xor_ln45_471_fu_13236_p2;
wire   [1:0] xor_ln45_436_fu_13248_p2;
wire   [1:0] xor_ln45_437_fu_13254_p2;
wire   [0:0] z1_170_fu_13273_p2;
wire   [0:0] z0_170_fu_13268_p2;
wire   [0:0] z2_168_fu_13278_p2;
wire   [0:0] xor_ln45_438_fu_13283_p2;
wire   [0:0] xor_ln45_439_fu_13289_p2;
wire   [0:0] z1_171_fu_13308_p2;
wire   [0:0] z0_172_fu_13303_p2;
wire   [0:0] z2_169_fu_13313_p2;
wire   [0:0] xor_ln45_440_fu_13318_p2;
wire   [0:0] xor_ln45_441_fu_13324_p2;
wire   [0:0] z1_173_fu_13343_p2;
wire   [0:0] z0_173_fu_13338_p2;
wire   [0:0] z2_170_fu_13348_p2;
wire   [0:0] a1_252_fu_13353_p2;
wire   [0:0] a0_278_fu_13359_p2;
wire   [0:0] xor_ln28_89_fu_13373_p2;
wire   [1:0] z1_172_fu_13330_p3;
wire   [1:0] z0_171_fu_13295_p3;
wire   [1:0] z2_225_fu_13365_p3;
wire   [1:0] tmp_88_fu_13379_p3;
wire   [1:0] xor_ln45_476_fu_13393_p2;
wire   [1:0] xor_ln45_475_fu_13387_p2;
wire   [1:0] a1_413_fu_13399_p2;
wire   [1:0] a0_279_fu_13405_p2;
wire   [0:0] a0_280_fu_13419_p1;
wire   [0:0] a1_254_fu_13423_p3;
wire   [0:0] xor_ln28_90_fu_13431_p2;
wire   [1:0] tmp_89_fu_13437_p3;
wire   [1:0] xor_ln28_91_fu_13445_p2;
wire   [3:0] z1_169_fu_13260_p3;
wire   [3:0] z0_165_fu_13109_p3;
wire   [3:0] z2_226_fu_13411_p3;
wire   [3:0] tmp_90_fu_13451_p3;
wire   [3:0] xor_ln45_480_fu_13465_p2;
wire   [3:0] xor_ln45_479_fu_13459_p2;
wire   [3:0] a1_414_fu_13471_p2;
wire   [3:0] a0_281_fu_13477_p2;
wire   [0:0] a0_283_fu_13505_p3;
wire   [0:0] a1_257_fu_13513_p3;
wire   [0:0] xor_ln28_92_fu_13521_p2;
wire   [1:0] a0_282_fu_13491_p1;
wire   [1:0] tmp_91_fu_13527_p3;
wire   [1:0] xor_ln28_93_fu_13535_p2;
wire   [1:0] a1_415_fu_13495_p4;
wire   [3:0] tmp_92_fu_13541_p3;
wire   [3:0] xor_ln28_94_fu_13549_p2;
wire   [7:0] z1_160_fu_12958_p3;
wire   [7:0] z0_147_fu_12433_p3;
wire   [7:0] z2_227_fu_13483_p3;
wire   [7:0] tmp_93_fu_13555_p3;
wire   [7:0] xor_ln45_484_fu_13569_p2;
wire   [7:0] xor_ln45_483_fu_13563_p2;
wire   [7:0] xor_ln45_348_fu_11904_p2;
wire   [7:0] xor_ln45_349_fu_11910_p2;
wire   [7:0] xor_ln45_454_fu_13575_p2;
wire   [7:0] xor_ln45_455_fu_13581_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_reset_idle_pp0;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        a0_288_reg_13599 <= a[32'd30];
        a0_288_reg_13599_pp0_iter1_reg <= a0_288_reg_13599;
        a0_329_reg_14028 <= a[32'd16];
        a0_329_reg_14028_pp0_iter1_reg <= a0_329_reg_14028;
        a0_330_reg_14046 <= a[32'd18];
        a0_330_reg_14046_pp0_iter1_reg <= a0_330_reg_14046;
        a0_331_reg_14057 <= a0_331_fu_4202_p2;
        a0_331_reg_14057_pp0_iter1_reg <= a0_331_reg_14057;
        a0_332_reg_14062 <= a[32'd20];
        a0_332_reg_14062_pp0_iter1_reg <= a0_332_reg_14062;
        a0_333_reg_14079 <= a[32'd22];
        a0_333_reg_14079_pp0_iter1_reg <= a0_333_reg_14079;
        a0_334_reg_14090 <= a0_334_fu_4286_p2;
        a0_334_reg_14090_pp0_iter1_reg <= a0_334_reg_14090;
        a0_335_reg_13615 <= a[32'd24];
        a0_335_reg_13615_pp0_iter1_reg <= a0_335_reg_13615;
        a0_336_reg_14105 <= a[32'd26];
        a0_336_reg_14105_pp0_iter1_reg <= a0_336_reg_14105;
        a0_337_reg_14116 <= a0_337_fu_4392_p2;
        a0_337_reg_14116_pp0_iter1_reg <= a0_337_reg_14116;
        a0_338_reg_14121 <= a[32'd28];
        a0_338_reg_14121_pp0_iter1_reg <= a0_338_reg_14121;
        a0_339_reg_13610 <= a0_339_fu_260_p2;
        a0_339_reg_13610_pp0_iter1_reg <= a0_339_reg_13610;
        a0_343_reg_14138 <= delta_fu_4668_p2[32'd14];
        a0_343_reg_14138_pp0_iter1_reg <= a0_343_reg_14138;
        a0_346_reg_14167 <= a0_346_fu_4922_p2;
        a0_348_reg_14197 <= a0_344_fu_4964_p2[32'd2];
        a0_352_reg_14268 <= a_170_fu_5142_p2[32'd2];
        a0_354_reg_14238 <= a0_340_fu_4704_p2[32'd4];
        a0_356_reg_14322 <= a0_340_fu_4704_p2[32'd6];
        a0_357_reg_14363 <= xor_ln71_3_fu_4686_p2[32'd8];
        a0_357_reg_14363_pp0_iter1_reg <= a0_357_reg_14363;
        a0_358_reg_14378 <= xor_ln71_3_fu_4686_p2[32'd10];
        a0_358_reg_14378_pp0_iter1_reg <= a0_358_reg_14378;
        a0_359_reg_14675 <= a0_359_fu_6635_p2;
        a0_360_reg_14159 <= delta_fu_4668_p2[32'd12];
        a0_360_reg_14159_pp0_iter1_reg <= a0_360_reg_14159;
        a0_361_reg_14151 <= a0_361_fu_4772_p2;
        a0_361_reg_14151_pp0_iter1_reg <= a0_361_reg_14151;
        a0_364_reg_14685 <= delta_1_fu_6731_p2[32'd6];
        a0_369_reg_14746 <= xor_ln71_4_fu_6737_p2[32'd4];
        a0_370_reg_14696 <= a0_370_fu_6785_p2;
        a0_377_reg_14784 <= a0_377_fu_7546_p2;
        a0_379_reg_14769 <= a0_379_fu_7516_p2;
        a1_261_reg_13605 <= a[32'd31];
        a1_261_reg_13605_pp0_iter1_reg <= a1_261_reg_13605;
        a1_307_reg_14036 <= a[32'd17];
        a1_307_reg_14036_pp0_iter1_reg <= a1_307_reg_14036;
        a1_308_reg_14052 <= a[32'd19];
        a1_308_reg_14052_pp0_iter1_reg <= a1_308_reg_14052;
        a1_309_reg_14069 <= a[32'd21];
        a1_309_reg_14069_pp0_iter1_reg <= a1_309_reg_14069;
        a1_310_reg_14085 <= a[32'd23];
        a1_310_reg_14085_pp0_iter1_reg <= a1_310_reg_14085;
        a1_311_reg_14095 <= a[32'd25];
        a1_311_reg_14095_pp0_iter1_reg <= a1_311_reg_14095;
        a1_312_reg_14111 <= a[32'd27];
        a1_312_reg_14111_pp0_iter1_reg <= a1_312_reg_14111;
        a1_313_reg_14128 <= a[32'd29];
        a1_313_reg_14128_pp0_iter1_reg <= a1_313_reg_14128;
        a1_318_reg_14145 <= delta_fu_4668_p2[32'd15];
        a1_318_reg_14145_pp0_iter1_reg <= a1_318_reg_14145;
        a1_321_reg_14175 <= a0_345_fu_4946_p2[32'd1];
        a1_322_reg_14212 <= a_161_fu_5072_p2[32'd1];
        a1_323_reg_14225 <= a0_344_fu_4964_p2[32'd3];
        a1_325_reg_14255 <= a0_349_fu_5172_p2[32'd1];
        a1_326_reg_14283 <= a_175_fu_5228_p2[32'd1];
        a1_327_reg_14296 <= a_170_fu_5142_p2[32'd3];
        a1_329_reg_14309 <= xor_ln68_3_fu_4710_p2[32'd5];
        a1_330_reg_14337 <= a_189_fu_5324_p2[32'd1];
        a1_331_reg_14350 <= a0_340_fu_4704_p2[32'd7];
        a1_333_reg_14371 <= xor_ln71_2_fu_4680_p2[32'd9];
        a1_333_reg_14371_pp0_iter1_reg <= a1_333_reg_14371;
        a1_334_reg_14385 <= xor_ln71_3_fu_4686_p2[32'd11];
        a1_334_reg_14385_pp0_iter1_reg <= a1_334_reg_14385;
        a1_335_reg_14397 <= xor_ln71_1_fu_4674_p2[32'd13];
        a1_335_reg_14397_pp0_iter1_reg <= a1_335_reg_14397;
        a1_337_reg_14691 <= delta_1_fu_6731_p2[32'd7];
        a1_342_reg_14752 <= xor_ln71_4_fu_6737_p2[32'd5];
        a1_348_reg_14777 <= a1_348_fu_7540_p2;
        a1_350_reg_14762 <= a1_350_fu_7510_p2;
        a_233_reg_14792 <= a_233_fu_7552_p2;
        a_241_reg_14804 <= a_241_fu_7572_p2;
        b0_11_reg_13668 <= b0_fu_484_p2[32'd4];
        b0_11_reg_13668_pp0_iter1_reg <= b0_11_reg_13668;
        b0_12_reg_13733 <= b0_12_fu_1352_p2;
        b0_12_reg_13733_pp0_iter1_reg <= b0_12_reg_13733;
        b0_13_reg_13728 <= b0_fu_484_p2[32'd6];
        b0_13_reg_13728_pp0_iter1_reg <= b0_13_reg_13728;
        b0_16_reg_13763 <= b0_16_fu_1802_p2;
        b0_16_reg_13763_pp0_iter1_reg <= b0_16_reg_13763;
        b0_17_reg_13783 <= b0_17_fu_1908_p2;
        b0_17_reg_13783_pp0_iter1_reg <= b0_17_reg_13783;
        b0_18_reg_13778 <= b0_14_fu_1740_p2[32'd2];
        b0_18_reg_13778_pp0_iter1_reg <= b0_18_reg_13778;
        b0_20_reg_13813 <= b0_20_fu_2178_p2;
        b0_20_reg_13813_pp0_iter1_reg <= b0_20_reg_13813;
        b0_21_reg_13833 <= b0_21_fu_2284_p2;
        b0_21_reg_13833_pp0_iter1_reg <= b0_21_reg_13833;
        b0_22_reg_13828 <= b_55_fu_2126_p2[32'd2];
        b0_22_reg_13828_pp0_iter1_reg <= b0_22_reg_13828;
        b0_24_reg_13808 <= b_41_fu_1712_p2[32'd4];
        b0_24_reg_13808_pp0_iter1_reg <= b0_24_reg_13808;
        b0_25_reg_13873 <= b0_25_fu_2588_p2;
        b0_25_reg_13873_pp0_iter1_reg <= b0_25_reg_13873;
        b0_26_reg_13868 <= b_41_fu_1712_p2[32'd6];
        b0_26_reg_13868_pp0_iter1_reg <= b0_26_reg_13868;
        b0_29_reg_13758 <= a0z1_fu_440_p2[32'd8];
        b0_29_reg_13758_pp0_iter1_reg <= b0_29_reg_13758;
        b0_30_reg_13913 <= b0_30_fu_3008_p2;
        b0_30_reg_13913_pp0_iter1_reg <= b0_30_reg_13913;
        b0_31_reg_13908 <= xor_ln70_3_fu_458_p2[32'd10];
        b0_31_reg_13908_pp0_iter1_reg <= b0_31_reg_13908;
        b0_33_reg_13943 <= b0_33_fu_3278_p2;
        b0_33_reg_13943_pp0_iter1_reg <= b0_33_reg_13943;
        b0_34_reg_13963 <= b0_34_fu_3384_p2;
        b0_34_reg_13963_pp0_iter1_reg <= b0_34_reg_13963;
        b0_35_reg_13958 <= b_95_fu_3226_p2[32'd2];
        b0_35_reg_13958_pp0_iter1_reg <= b0_35_reg_13958;
        b0_37_reg_13938 <= a0z1_fu_440_p2[32'd12];
        b0_37_reg_13938_pp0_iter1_reg <= b0_37_reg_13938;
        b0_38_reg_14003 <= b0_38_fu_3688_p2;
        b0_38_reg_14003_pp0_iter1_reg <= b0_38_reg_14003;
        b0_39_reg_13998 <= a0z1_fu_440_p2[32'd14];
        b0_39_reg_13998_pp0_iter1_reg <= b0_39_reg_13998;
        b0_3_reg_13623 <= b0_3_fu_566_p2;
        b0_3_reg_13623_pp0_iter1_reg <= b0_3_reg_13623;
        b0_42_reg_14181 <= b0_42_fu_5050_p2;
        b0_42_reg_14181_pp0_iter1_reg <= b0_42_reg_14181;
        b0_43_reg_14610 <= b0_43_fu_6014_p2;
        b0_44_reg_14204 <= b0_40_fu_5000_p2[32'd2];
        b0_44_reg_14204_pp0_iter1_reg <= b0_44_reg_14204;
        b0_46_reg_14625 <= b0_46_fu_6156_p2;
        b0_47_reg_14635 <= b0_47_fu_6211_p2;
        b0_48_reg_14275 <= b_135_fu_5166_p2[32'd2];
        b0_48_reg_14275_pp0_iter1_reg <= b0_48_reg_14275;
        b0_4_reg_13643 <= b0_4_fu_672_p2;
        b0_4_reg_13643_pp0_iter1_reg <= b0_4_reg_13643;
        b0_50_reg_14246 <= a0z1_1_fu_4978_p2[32'd4];
        b0_50_reg_14246_pp0_iter1_reg <= b0_50_reg_14246;
        b0_51_reg_14655 <= b0_51_fu_6396_p2;
        b0_52_reg_14329 <= a0z1_1_fu_4978_p2[32'd6];
        b0_52_reg_14329_pp0_iter1_reg <= b0_52_reg_14329;
        b0_54_reg_14701 <= b0_54_fu_6912_p2;
        b0_55_reg_14721 <= b0_55_fu_7018_p2;
        b0_56_reg_14716 <= a0z1_2_fu_6872_p2[32'd2];
        b0_5_reg_13638 <= b0_1_fu_516_p2[32'd2];
        b0_5_reg_13638_pp0_iter1_reg <= b0_5_reg_13638;
        b0_64_reg_14423 <= b_208_fu_5460_p2[32'd2];
        b0_64_reg_14423_pp0_iter1_reg <= b0_64_reg_14423;
        b0_72_reg_14460 <= b_248_fu_5578_p2[32'd2];
        b0_72_reg_14460_pp0_iter1_reg <= b0_72_reg_14460;
        b0_79_reg_14491 <= b0_75_fu_5674_p2[32'd2];
        b0_79_reg_14491_pp0_iter1_reg <= b0_79_reg_14491;
        b0_7_reg_13673 <= b0_7_fu_942_p2;
        b0_7_reg_13673_pp0_iter1_reg <= b0_7_reg_13673;
        b0_83_reg_14524 <= b_288_fu_5762_p2[32'd2];
        b0_83_reg_14524_pp0_iter1_reg <= b0_83_reg_14524;
        b0_85_reg_14510 <= b_274_fu_5662_p2[32'd4];
        b0_85_reg_14510_pp0_iter1_reg <= b0_85_reg_14510;
        b0_87_reg_14549 <= b_274_fu_5662_p2[32'd6];
        b0_87_reg_14549_pp0_iter1_reg <= b0_87_reg_14549;
        b0_8_reg_13693 <= b0_8_fu_1048_p2;
        b0_8_reg_13693_pp0_iter1_reg <= b0_8_reg_13693;
        b0_93_reg_14580 <= b_328_fu_5894_p2[32'd2];
        b0_93_reg_14580_pp0_iter1_reg <= b0_93_reg_14580;
        b0_9_reg_13688 <= b_15_fu_890_p2[32'd2];
        b0_9_reg_13688_pp0_iter1_reg <= b0_9_reg_13688;
        b1_100_reg_13648 <= b_7_fu_652_p2[32'd1];
        b1_100_reg_13648_pp0_iter1_reg <= b1_100_reg_13648;
        b1_101_reg_13658 <= b0_1_fu_516_p2[32'd3];
        b1_101_reg_13658_pp0_iter1_reg <= b1_101_reg_13658;
        b1_103_reg_13678 <= b0_6_fu_912_p2[32'd1];
        b1_103_reg_13678_pp0_iter1_reg <= b1_103_reg_13678;
        b1_104_reg_13698 <= b_20_fu_1028_p2[32'd1];
        b1_104_reg_13698_pp0_iter1_reg <= b1_104_reg_13698;
        b1_105_reg_13708 <= b_15_fu_890_p2[32'd3];
        b1_105_reg_13708_pp0_iter1_reg <= b1_105_reg_13708;
        b1_107_reg_13718 <= xor_ln40_1_fu_490_p2[32'd5];
        b1_107_reg_13718_pp0_iter1_reg <= b1_107_reg_13718;
        b1_108_reg_13738 <= b_33_fu_1332_p2[32'd1];
        b1_108_reg_13738_pp0_iter1_reg <= b1_108_reg_13738;
        b1_109_reg_13748 <= b0_fu_484_p2[32'd7];
        b1_109_reg_13748_pp0_iter1_reg <= b1_109_reg_13748;
        b1_112_reg_13768 <= b0_15_fu_1772_p2[32'd1];
        b1_112_reg_13768_pp0_iter1_reg <= b1_112_reg_13768;
        b1_113_reg_13788 <= b_47_fu_1888_p2[32'd1];
        b1_113_reg_13788_pp0_iter1_reg <= b1_113_reg_13788;
        b1_114_reg_13798 <= b0_14_fu_1740_p2[32'd3];
        b1_114_reg_13798_pp0_iter1_reg <= b1_114_reg_13798;
        b1_116_reg_13818 <= b0_19_fu_2148_p2[32'd1];
        b1_116_reg_13818_pp0_iter1_reg <= b1_116_reg_13818;
        b1_117_reg_13838 <= b_60_fu_2264_p2[32'd1];
        b1_117_reg_13838_pp0_iter1_reg <= b1_117_reg_13838;
        b1_118_reg_13848 <= b_55_fu_2126_p2[32'd3];
        b1_118_reg_13848_pp0_iter1_reg <= b1_118_reg_13848;
        b1_120_reg_13858 <= xor_ln33_fu_1718_p2[32'd5];
        b1_120_reg_13858_pp0_iter1_reg <= b1_120_reg_13858;
        b1_121_reg_13878 <= b_73_fu_2568_p2[32'd1];
        b1_121_reg_13878_pp0_iter1_reg <= b1_121_reg_13878;
        b1_122_reg_13888 <= b_41_fu_1712_p2[32'd7];
        b1_122_reg_13888_pp0_iter1_reg <= b1_122_reg_13888;
        b1_125_reg_13898 <= xor_ln70_2_fu_452_p2[32'd9];
        b1_125_reg_13898_pp0_iter1_reg <= b1_125_reg_13898;
        b1_126_reg_13918 <= b_87_fu_2988_p2[32'd1];
        b1_126_reg_13918_pp0_iter1_reg <= b1_126_reg_13918;
        b1_127_reg_13928 <= xor_ln70_3_fu_458_p2[32'd11];
        b1_127_reg_13928_pp0_iter1_reg <= b1_127_reg_13928;
        b1_129_reg_13948 <= b0_32_fu_3248_p2[32'd1];
        b1_129_reg_13948_pp0_iter1_reg <= b1_129_reg_13948;
        b1_130_reg_13968 <= b_100_fu_3364_p2[32'd1];
        b1_130_reg_13968_pp0_iter1_reg <= b1_130_reg_13968;
        b1_131_reg_13978 <= b_95_fu_3226_p2[32'd3];
        b1_131_reg_13978_pp0_iter1_reg <= b1_131_reg_13978;
        b1_133_reg_13988 <= xor_ln70_1_fu_446_p2[32'd13];
        b1_133_reg_13988_pp0_iter1_reg <= b1_133_reg_13988;
        b1_134_reg_14008 <= b_113_fu_3668_p2[32'd1];
        b1_134_reg_14008_pp0_iter1_reg <= b1_134_reg_14008;
        b1_135_reg_14018 <= a0z1_fu_440_p2[32'd15];
        b1_135_reg_14018_pp0_iter1_reg <= b1_135_reg_14018;
        b1_138_reg_14190 <= b0_41_fu_5026_p2[32'd1];
        b1_138_reg_14190_pp0_iter1_reg <= b1_138_reg_14190;
        b1_139_reg_14218 <= b_127_fu_5086_p2[32'd1];
        b1_139_reg_14218_pp0_iter1_reg <= b1_139_reg_14218;
        b1_140_reg_14231 <= b0_40_fu_5000_p2[32'd3];
        b1_140_reg_14231_pp0_iter1_reg <= b1_140_reg_14231;
        b1_142_reg_14261 <= b0_45_fu_5188_p2[32'd1];
        b1_142_reg_14261_pp0_iter1_reg <= b1_142_reg_14261;
        b1_143_reg_14289 <= b_140_fu_5242_p2[32'd1];
        b1_143_reg_14289_pp0_iter1_reg <= b1_143_reg_14289;
        b1_144_reg_14302 <= b_135_fu_5166_p2[32'd3];
        b1_144_reg_14302_pp0_iter1_reg <= b1_144_reg_14302;
        b1_146_reg_14315 <= xor_ln70_27_fu_4984_p2[32'd5];
        b1_146_reg_14315_pp0_iter1_reg <= b1_146_reg_14315;
        b1_147_reg_14343 <= b_153_fu_5338_p2[32'd1];
        b1_147_reg_14343_pp0_iter1_reg <= b1_147_reg_14343;
        b1_148_reg_14356 <= a0z1_1_fu_4978_p2[32'd7];
        b1_148_reg_14356_pp0_iter1_reg <= b1_148_reg_14356;
        b1_150_reg_14706 <= b0_53_fu_6888_p2[32'd1];
        b1_151_reg_14726 <= b_166_fu_6998_p2[32'd1];
        b1_152_reg_14736 <= a0z1_2_fu_6872_p2[32'd3];
        b1_154_reg_14798 <= b_187_fu_7558_p2[32'd1];
        b1_156_reg_14411 <= b_200_fu_5446_p2[32'd1];
        b1_156_reg_14411_pp0_iter1_reg <= b1_156_reg_14411;
        b1_158_reg_14417 <= b0_61_fu_5466_p2[32'd1];
        b1_158_reg_14417_pp0_iter1_reg <= b1_158_reg_14417;
        b1_159_reg_14430 <= b_213_fu_5498_p2[32'd1];
        b1_159_reg_14430_pp0_iter1_reg <= b1_159_reg_14430;
        b1_160_reg_14436 <= b_208_fu_5460_p2[32'd3];
        b1_160_reg_14436_pp0_iter1_reg <= b1_160_reg_14436;
        b1_161_reg_14442 <= b_226_fu_5520_p2[32'd1];
        b1_161_reg_14442_pp0_iter1_reg <= b1_161_reg_14442;
        b1_164_reg_14448 <= b_240_fu_5554_p2[32'd1];
        b1_164_reg_14448_pp0_iter1_reg <= b1_164_reg_14448;
        b1_166_reg_14454 <= b0_69_fu_5584_p2[32'd1];
        b1_166_reg_14454_pp0_iter1_reg <= b1_166_reg_14454;
        b1_167_reg_14467 <= b_253_fu_5616_p2[32'd1];
        b1_167_reg_14467_pp0_iter1_reg <= b1_167_reg_14467;
        b1_168_reg_14473 <= b_248_fu_5578_p2[32'd3];
        b1_168_reg_14473_pp0_iter1_reg <= b1_168_reg_14473;
        b1_170_reg_14479 <= b_266_fu_5648_p2[32'd1];
        b1_170_reg_14479_pp0_iter1_reg <= b1_170_reg_14479;
        b1_173_reg_14485 <= b0_76_fu_5690_p2[32'd1];
        b1_173_reg_14485_pp0_iter1_reg <= b1_173_reg_14485;
        b1_174_reg_14498 <= b_280_fu_5722_p2[32'd1];
        b1_174_reg_14498_pp0_iter1_reg <= b1_174_reg_14498;
        b1_175_reg_14504 <= b0_75_fu_5674_p2[32'd3];
        b1_175_reg_14504_pp0_iter1_reg <= b1_175_reg_14504;
        b1_177_reg_14518 <= b0_80_fu_5768_p2[32'd1];
        b1_177_reg_14518_pp0_iter1_reg <= b1_177_reg_14518;
        b1_178_reg_14531 <= b_293_fu_5800_p2[32'd1];
        b1_178_reg_14531_pp0_iter1_reg <= b1_178_reg_14531;
        b1_179_reg_14537 <= b_288_fu_5762_p2[32'd3];
        b1_179_reg_14537_pp0_iter1_reg <= b1_179_reg_14537;
        b1_181_reg_14543 <= xor_ln33_1_fu_5668_p2[32'd5];
        b1_181_reg_14543_pp0_iter1_reg <= b1_181_reg_14543;
        b1_182_reg_14556 <= b_306_fu_5848_p2[32'd1];
        b1_182_reg_14556_pp0_iter1_reg <= b1_182_reg_14556;
        b1_183_reg_14562 <= b_274_fu_5662_p2[32'd7];
        b1_183_reg_14562_pp0_iter1_reg <= b1_183_reg_14562;
        b1_185_reg_14568 <= b_320_fu_5880_p2[32'd1];
        b1_185_reg_14568_pp0_iter1_reg <= b1_185_reg_14568;
        b1_187_reg_14574 <= b0_90_fu_5900_p2[32'd1];
        b1_187_reg_14574_pp0_iter1_reg <= b1_187_reg_14574;
        b1_188_reg_14587 <= b_333_fu_5932_p2[32'd1];
        b1_188_reg_14587_pp0_iter1_reg <= b1_188_reg_14587;
        b1_189_reg_14593 <= b_328_fu_5894_p2[32'd3];
        b1_189_reg_14593_pp0_iter1_reg <= b1_189_reg_14593;
        b1_190_reg_14599 <= b_346_fu_5954_p2[32'd1];
        b1_190_reg_14599_pp0_iter1_reg <= b1_190_reg_14599;
        b1_99_reg_13628 <= b0_2_fu_542_p2[32'd1];
        b1_99_reg_13628_pp0_iter1_reg <= b1_99_reg_13628;
        b_102_reg_13973 <= b_102_fu_3410_p2;
        b_102_reg_13973_pp0_iter1_reg <= b_102_reg_13973;
        b_106_reg_13983 <= b_106_fu_3476_p2;
        b_106_reg_13983_pp0_iter1_reg <= b_106_reg_13983;
        b_111_reg_13993 <= b_111_fu_3608_p2;
        b_111_reg_13993_pp0_iter1_reg <= b_111_reg_13993;
        b_115_reg_14013 <= b_115_fu_3714_p2;
        b_115_reg_14013_pp0_iter1_reg <= b_115_reg_14013;
        b_119_reg_14023 <= b_119_fu_3780_p2;
        b_119_reg_14023_pp0_iter1_reg <= b_119_reg_14023;
        b_125_reg_14605 <= b_125_fu_5976_p2;
        b_129_reg_14615 <= b_129_fu_6029_p2;
        b_133_reg_14620 <= b_133_fu_6072_p2;
        b_138_reg_14630 <= b_138_fu_6171_p2;
        b_13_reg_13663 <= b_13_fu_764_p2;
        b_13_reg_13663_pp0_iter1_reg <= b_13_reg_13663;
        b_142_reg_14640 <= b_142_fu_6227_p2;
        b_146_reg_14645 <= b_146_fu_6270_p2;
        b_151_reg_14650 <= b_151_fu_6358_p2;
        b_155_reg_14660 <= b_155_fu_6411_p2;
        b_159_reg_14665 <= b_159_fu_6454_p2;
        b_164_reg_14711 <= b_164_fu_6938_p2;
        b_168_reg_14731 <= b_168_fu_7044_p2;
        b_172_reg_14741 <= b_172_fu_7110_p2;
        b_185_reg_14757 <= b_185_fu_7222_p2;
        b_18_reg_13683 <= b_18_fu_968_p2;
        b_18_reg_13683_pp0_iter1_reg <= b_18_reg_13683;
        b_198_reg_14670 <= b_198_fu_6624_p2;
        b_224_reg_14680 <= b_224_fu_6659_p2;
        b_22_reg_13703 <= b_22_fu_1074_p2;
        b_22_reg_13703_pp0_iter1_reg <= b_22_reg_13703;
        b_238_reg_14041 <= b_238_fu_4172_p2;
        b_238_reg_14041_pp0_iter1_reg <= b_238_reg_14041;
        b_264_reg_14074 <= b_264_fu_4256_p2;
        b_264_reg_14074_pp0_iter1_reg <= b_264_reg_14074;
        b_26_reg_13713 <= b_26_fu_1140_p2;
        b_26_reg_13713_pp0_iter1_reg <= b_26_reg_13713;
        b_318_reg_14100 <= b_318_fu_4362_p2;
        b_318_reg_14100_pp0_iter1_reg <= b_318_reg_14100;
        b_31_reg_13723 <= b_31_fu_1272_p2;
        b_31_reg_13723_pp0_iter1_reg <= b_31_reg_13723;
        b_344_reg_14133 <= b_344_fu_4446_p2;
        b_344_reg_14133_pp0_iter1_reg <= b_344_reg_14133;
        b_35_reg_13743 <= b_35_fu_1378_p2;
        b_35_reg_13743_pp0_iter1_reg <= b_35_reg_13743;
        b_39_reg_13753 <= b_39_fu_1444_p2;
        b_39_reg_13753_pp0_iter1_reg <= b_39_reg_13753;
        b_45_reg_13773 <= b_45_fu_1828_p2;
        b_45_reg_13773_pp0_iter1_reg <= b_45_reg_13773;
        b_49_reg_13793 <= b_49_fu_1934_p2;
        b_49_reg_13793_pp0_iter1_reg <= b_49_reg_13793;
        b_53_reg_13803 <= b_53_fu_2000_p2;
        b_53_reg_13803_pp0_iter1_reg <= b_53_reg_13803;
        b_58_reg_13823 <= b_58_fu_2204_p2;
        b_58_reg_13823_pp0_iter1_reg <= b_58_reg_13823;
        b_5_reg_13633 <= b_5_fu_592_p2;
        b_5_reg_13633_pp0_iter1_reg <= b_5_reg_13633;
        b_62_reg_13843 <= b_62_fu_2310_p2;
        b_62_reg_13843_pp0_iter1_reg <= b_62_reg_13843;
        b_66_reg_13853 <= b_66_fu_2376_p2;
        b_66_reg_13853_pp0_iter1_reg <= b_66_reg_13853;
        b_71_reg_13863 <= b_71_fu_2508_p2;
        b_71_reg_13863_pp0_iter1_reg <= b_71_reg_13863;
        b_75_reg_13883 <= b_75_fu_2614_p2;
        b_75_reg_13883_pp0_iter1_reg <= b_75_reg_13883;
        b_79_reg_13893 <= b_79_fu_2680_p2;
        b_79_reg_13893_pp0_iter1_reg <= b_79_reg_13893;
        b_85_reg_13903 <= b_85_fu_2928_p2;
        b_85_reg_13903_pp0_iter1_reg <= b_85_reg_13903;
        b_89_reg_13923 <= b_89_fu_3034_p2;
        b_89_reg_13923_pp0_iter1_reg <= b_89_reg_13923;
        b_93_reg_13933 <= b_93_fu_3100_p2;
        b_93_reg_13933_pp0_iter1_reg <= b_93_reg_13933;
        b_98_reg_13953 <= b_98_fu_3304_p2;
        b_98_reg_13953_pp0_iter1_reg <= b_98_reg_13953;
        b_9_reg_13653 <= b_9_fu_698_p2;
        b_9_reg_13653_pp0_iter1_reg <= b_9_reg_13653;
        tmp_256_reg_14392 <= tmp_256_fu_5408_p4;
        tmp_258_reg_14404 <= tmp_258_fu_5426_p4;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

assign ap_reset_idle_pp0 = 1'b0;

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign a0_111_fu_6092_p2 = (z2_42_fu_6082_p2 ^ z0_43_fu_6064_p2);

assign a0_117_fu_6290_p2 = (z2_46_fu_6280_p2 ^ z0_48_fu_6262_p2);

assign a0_128_fu_6474_p2 = (z2_50_fu_6464_p2 ^ z0_52_fu_6446_p2);

assign a0_129_fu_6520_p2 = (z2_189_fu_6480_p3 ^ z0_50_fu_6384_p3);

assign a0_130_fu_6534_p1 = a1_332_fu_6514_p2[0:0];

assign a0_138_fu_6676_p2 = (a1_sqr_32_fu_6670_p3 ^ a0_sqr_20_fu_6663_p3);

assign a0_150_fu_7134_p2 = (z2_55_fu_7122_p2 ^ z0_56_fu_7098_p2);

assign a0_167_fu_7710_p2 = (z2_62_fu_7700_p2 ^ z0_63_fu_7692_p2);

assign a0_16_fu_1164_p2 = (z2_6_fu_1152_p2 ^ z0_8_fu_1128_p2);

assign a0_170_fu_7847_p2 = (z2_66_fu_7837_p2 ^ z0_67_fu_7829_p2);

assign a0_190_fu_8069_p2 = (z2_70_fu_8058_p2 ^ z0_71_fu_8042_p2);

assign a0_195_fu_8342_p2 = (z2_74_fu_8331_p2 ^ z0_76_fu_8310_p2);

assign a0_200_fu_8562_p2 = (z2_78_fu_8551_p2 ^ z0_80_fu_8535_p2);

assign a0_201_fu_8608_p2 = (z2_196_fu_8568_p3 ^ z0_78_fu_8443_p3);

assign a0_202_fu_8622_p1 = a1_364_fu_8602_p2[0:0];

assign a0_203_fu_8789_p2 = (z2_83_fu_8778_p2 ^ z0_84_fu_8768_p2);

assign a0_204_fu_8940_p2 = (z2_87_fu_8929_p2 ^ z0_89_fu_8919_p2);

assign a0_205_fu_9091_p2 = (z2_91_fu_9080_p2 ^ z0_93_fu_9070_p2);

assign a0_206_fu_9137_p2 = (z2_200_fu_9097_p3 ^ z0_91_fu_9027_p3);

assign a0_207_fu_9151_p1 = a1_365_fu_9131_p2[0:0];

assign a0_214_fu_9455_p2 = (z2_96_fu_9444_p2 ^ z0_97_fu_9428_p2);

assign a0_219_fu_9726_p2 = (z2_100_fu_9715_p2 ^ z0_102_fu_9694_p2);

assign a0_224_fu_9960_p2 = (z2_104_fu_9949_p2 ^ z0_106_fu_9933_p2);

assign a0_225_fu_10006_p2 = (z2_204_fu_9966_p3 ^ z0_104_fu_9837_p3);

assign a0_226_fu_10020_p1 = a1_380_fu_10000_p2[0:0];

assign a0_232_fu_10343_p2 = (z2_109_fu_10332_p2 ^ z0_111_fu_10311_p2);

assign a0_237_fu_10631_p2 = (z2_113_fu_10620_p2 ^ z0_116_fu_10599_p2);

assign a0_23_fu_1468_p2 = (z2_10_fu_1456_p2 ^ z0_12_fu_1432_p2);

assign a0_242_fu_10875_p2 = (z2_117_fu_10864_p2 ^ z0_120_fu_10843_p2);

assign a0_243_fu_10921_p2 = (z2_208_fu_10881_p3 ^ z0_118_fu_10747_p3);

assign a0_244_fu_10935_p1 = a1_394_fu_10915_p2[0:0];

assign a0_24_fu_1514_p2 = (z2_176_fu_1474_p3 ^ z0_10_fu_1302_p3);

assign a0_250_fu_11181_p2 = (z2_122_fu_11170_p2 ^ z0_124_fu_11154_p2);

assign a0_255_fu_11454_p2 = (z2_126_fu_11443_p2 ^ z0_129_fu_11422_p2);

assign a0_25_fu_1528_p1 = a1_276_fu_1508_p2[0:0];

assign a0_260_fu_11688_p2 = (z2_130_fu_11677_p2 ^ z0_133_fu_11661_p2);

assign a0_261_fu_11734_p2 = (z2_212_fu_11694_p3 ^ z0_131_fu_11565_p3);

assign a0_262_fu_11748_p1 = a1_408_fu_11728_p2[0:0];

assign a0_263_fu_11806_p2 = (z2_213_fu_11740_p3 ^ z0_125_fu_11233_p3);

assign a0_264_fu_11820_p1 = a1_409_fu_11800_p2[1:0];

assign a0_265_fu_11834_p3 = a1_409_fu_11800_p2[32'd2];

assign a0_266_fu_12007_p2 = (z2_136_fu_11996_p2 ^ z0_137_fu_11986_p2);

assign a0_267_fu_12158_p2 = (z2_140_fu_12147_p2 ^ z0_142_fu_12137_p2);

assign a0_268_fu_12309_p2 = (z2_144_fu_12298_p2 ^ z0_146_fu_12288_p2);

assign a0_269_fu_12355_p2 = (z2_217_fu_12315_p3 ^ z0_144_fu_12245_p3);

assign a0_270_fu_12369_p1 = a1_411_fu_12349_p2[0:0];

assign a0_271_fu_12532_p2 = (z2_149_fu_12521_p2 ^ z0_151_fu_12511_p2);

assign a0_272_fu_12683_p2 = (z2_153_fu_12672_p2 ^ z0_156_fu_12662_p2);

assign a0_273_fu_12834_p2 = (z2_157_fu_12823_p2 ^ z0_160_fu_12813_p2);

assign a0_274_fu_12880_p2 = (z2_221_fu_12840_p3 ^ z0_158_fu_12770_p3);

assign a0_275_fu_12894_p1 = a1_412_fu_12874_p2[0:0];

assign a0_276_fu_13057_p2 = (z2_162_fu_13046_p2 ^ z0_164_fu_13036_p2);

assign a0_277_fu_13208_p2 = (z2_166_fu_13197_p2 ^ z0_169_fu_13187_p2);

assign a0_278_fu_13359_p2 = (z2_170_fu_13348_p2 ^ z0_173_fu_13338_p2);

assign a0_279_fu_13405_p2 = (z2_225_fu_13365_p3 ^ z0_171_fu_13295_p3);

assign a0_280_fu_13419_p1 = a1_413_fu_13399_p2[0:0];

assign a0_281_fu_13477_p2 = (z2_226_fu_13411_p3 ^ z0_165_fu_13109_p3);

assign a0_282_fu_13491_p1 = a1_414_fu_13471_p2[1:0];

assign a0_283_fu_13505_p3 = a1_414_fu_13471_p2[32'd2];

assign a0_284_fu_168_p1 = a[15:0];

assign a0_285_fu_184_p4 = {{a[23:16]}};

assign a0_286_fu_204_p4 = {{a[27:24]}};

assign a0_287_fu_224_p4 = {{a[29:28]}};

assign a0_288_fu_244_p3 = a[32'd30];

assign a0_289_fu_408_p1 = a[7:0];

assign a0_290_fu_404_p1 = a[3:0];

assign a0_291_fu_400_p1 = a[1:0];

assign a0_292_fu_396_p1 = a[0:0];

assign a0_293_fu_658_p2 = (a0_294_fu_630_p3 ^ a0_292_fu_396_p1);

assign a0_294_fu_630_p3 = a[32'd2];

assign a0_295_fu_896_p2 = (a0_299_fu_856_p4 ^ a0_291_fu_400_p1);

assign a0_296_fu_928_p2 = (a0_300_fu_848_p3 ^ a0_292_fu_396_p1);

assign a0_297_fu_1034_p2 = (a0_298_fu_1006_p3 ^ a0_296_fu_928_p2);

assign a0_298_fu_1006_p3 = a_20_fu_866_p2[32'd2];

assign a0_299_fu_856_p4 = {{a[5:4]}};

assign a0_300_fu_848_p3 = a[32'd4];

assign a0_301_fu_1338_p2 = (a0_302_fu_1310_p3 ^ a0_300_fu_848_p3);

assign a0_302_fu_1310_p3 = a[32'd6];

assign a0_303_fu_1724_p2 = (a0_316_fu_1642_p4 ^ a0_290_fu_404_p1);

assign a0_304_fu_1756_p2 = (a0_317_fu_1632_p4 ^ a0_291_fu_400_p1);

assign a0_305_fu_1788_p2 = (a0_318_fu_1624_p3 ^ a0_292_fu_396_p1);

assign a0_306_fu_1894_p2 = (a0_307_fu_1866_p3 ^ a0_305_fu_1788_p2);

assign a0_307_fu_1866_p3 = a0_303_fu_1724_p2[32'd2];

assign a0_308_fu_2132_p2 = (a0_312_fu_2092_p4 ^ a0_304_fu_1756_p2);

assign a0_309_fu_2164_p2 = (a0_313_fu_2084_p3 ^ a0_305_fu_1788_p2);

assign a0_310_fu_2270_p2 = (a0_311_fu_2242_p3 ^ a0_309_fu_2164_p2);

assign a0_311_fu_2242_p3 = a_65_fu_2102_p2[32'd2];

assign a0_312_fu_2092_p4 = {{a_50_fu_1662_p2[5:4]}};

assign a0_313_fu_2084_p3 = a_50_fu_1662_p2[32'd4];

assign a0_314_fu_2574_p2 = (a0_315_fu_2546_p3 ^ a0_313_fu_2084_p3);

assign a0_315_fu_2546_p3 = a_50_fu_1662_p2[32'd6];

assign a0_316_fu_1642_p4 = {{a[11:8]}};

assign a0_317_fu_1632_p4 = {{a[9:8]}};

assign a0_318_fu_1624_p3 = a[32'd8];

assign a0_319_fu_2994_p2 = (a0_320_fu_2966_p3 ^ a0_318_fu_1624_p3);

assign a0_320_fu_2966_p3 = a[32'd10];

assign a0_321_fu_3232_p2 = (a0_325_fu_3192_p4 ^ a0_317_fu_1632_p4);

assign a0_322_fu_3264_p2 = (a0_326_fu_3184_p3 ^ a0_318_fu_1624_p3);

assign a0_323_fu_3370_p2 = (a0_324_fu_3342_p3 ^ a0_322_fu_3264_p2);

assign a0_324_fu_3342_p3 = a_110_fu_3202_p2[32'd2];

assign a0_325_fu_3192_p4 = {{a[13:12]}};

assign a0_326_fu_3184_p3 = a[32'd12];

assign a0_327_fu_3674_p2 = (a0_328_fu_3646_p3 ^ a0_326_fu_3184_p3);

assign a0_328_fu_3646_p3 = a[32'd14];

assign a0_329_fu_4156_p3 = a[32'd16];

assign a0_330_fu_4186_p3 = a[32'd18];

assign a0_331_fu_4202_p2 = (a1_308_fu_4194_p3 ^ a0_330_fu_4186_p3);

assign a0_332_fu_4240_p3 = a[32'd20];

assign a0_333_fu_4270_p3 = a[32'd22];

assign a0_334_fu_4286_p2 = (a1_310_fu_4278_p3 ^ a0_333_fu_4270_p3);

assign a0_335_fu_362_p3 = a[32'd24];

assign a0_336_fu_4376_p3 = a[32'd26];

assign a0_337_fu_4392_p2 = (a1_312_fu_4384_p3 ^ a0_336_fu_4376_p3);

assign a0_338_fu_4430_p3 = a[32'd28];

assign a0_339_fu_260_p2 = (a1_261_fu_252_p3 ^ a0_288_fu_244_p3);

assign a0_340_fu_4704_p2 = (xor_ln59_13_fu_4590_p2 ^ xor_ln45_105_fu_4124_p2);

assign a0_341_fu_4716_p4 = {{xor_ln71_3_fu_4686_p2[11:8]}};

assign a0_342_fu_4736_p4 = {{delta_fu_4668_p2[13:12]}};

assign a0_343_fu_4756_p3 = delta_fu_4668_p2[32'd14];

assign a0_344_fu_4964_p2 = (xor_ln70_24_fu_4958_p2 ^ xor_ln70_23_fu_4952_p2);

assign a0_345_fu_4946_p2 = (xor_ln70_21_fu_4940_p2 ^ xor_ln70_20_fu_4934_p2);

assign a0_346_fu_4922_p2 = (xor_ln70_9_fu_4874_p2 ^ xor_ln70_16_fu_4916_p2);

assign a0_347_fu_6010_p2 = (a0_348_reg_14197 ^ a0_346_reg_14167);

assign a0_349_fu_5172_p2 = (a0_353_fu_5132_p4 ^ a0_345_fu_4946_p2);

assign a0_350_fu_6152_p2 = (a0_354_reg_14238 ^ a0_346_reg_14167);

assign a0_351_fu_6206_p2 = (a0_352_reg_14268 ^ a0_350_fu_6152_p2);

assign a0_353_fu_5132_p4 = {{a0_340_fu_4704_p2[5:4]}};

assign a0_355_fu_6392_p2 = (a0_356_reg_14322 ^ a0_354_reg_14238);

assign a0_359_fu_6635_p2 = (a1_334_reg_14385 ^ a0_358_reg_14378);

assign a0_360_fu_4816_p3 = delta_fu_4668_p2[32'd12];

assign a0_361_fu_4772_p2 = (a1_318_fu_4764_p3 ^ a0_343_fu_4756_p3);

assign a0_362_fu_6743_p2 = (xor_ln59_19_fu_6701_p2 ^ xor_ln45_139_fu_6604_p2);

assign a0_363_fu_6749_p4 = {{xor_ln71_4_fu_6737_p2[5:4]}};

assign a0_364_fu_6769_p3 = delta_1_fu_6731_p2[32'd6];

assign a0_365_fu_6866_p2 = (xor_ln70_36_fu_6860_p2 ^ xor_ln70_35_fu_6854_p2);

assign a0_366_fu_6848_p2 = (xor_ln70_33_fu_6842_p2 ^ xor_ln70_30_fu_6824_p2);

assign a0_367_fu_7004_p2 = (a0_368_fu_6976_p3 ^ a0_366_fu_6848_p2);

assign a0_368_fu_6976_p3 = a0_362_fu_6743_p2[32'd2];

assign a0_369_fu_7206_p3 = xor_ln71_4_fu_6737_p2[32'd4];

assign a0_36_fu_2024_p2 = (z2_15_fu_2012_p2 ^ z0_17_fu_1988_p2);

assign a0_370_fu_6785_p2 = (a1_337_fu_6777_p3 ^ a0_364_fu_6769_p3);

assign a0_371_fu_7314_p2 = (xor_ln59_21_fu_7244_p2 ^ xor_ln45_149_fu_7186_p2);

assign a0_372_fu_7320_p3 = xor_ln36_fu_7290_p2[32'd2];

assign a0_373_fu_7308_p2 = (xor_ln36_2_fu_7302_p2 ^ xor_ln36_1_fu_7296_p2);

assign a0_374_fu_7442_p2 = (xor_ln45_151_fu_7414_p2 ^ b_181_fu_7336_p2);

assign a0_375_fu_7480_p2 = (delta_4_fu_7468_p2 & a0z1_4_fu_7456_p2);

assign a0_376_fu_7578_p3 = {{a1_348_reg_14777}, {a0_377_reg_14784}};

assign a0_377_fu_7546_p2 = (z2_59_fu_7534_p2 ^ z0_59_fu_7522_p2);

assign a0_378_fu_7628_p2 = (a0_379_reg_14769 ^ a0_377_reg_14784);

assign a0_379_fu_7516_p2 = (z2_58_fu_7504_p2 ^ z0_58_fu_7486_p2);

assign a0_380_fu_7899_p3 = {{a1_352_fu_7887_p2}, {a0_381_fu_7875_p2}};

assign a0_381_fu_7875_p2 = (z2_193_fu_7853_p3 ^ z0_65_fu_7786_p3);

assign a0_382_fu_7893_p2 = (xor_ln45_167_fu_7780_p2 ^ a0_170_fu_7847_p2);

assign a0_383_fu_7968_p2 = (a0_384_fu_7964_p1 ^ a0_382_fu_7893_p2);

assign a0_384_fu_7964_p1 = a1_352_fu_7887_p2[0:0];

assign a0_385_fu_8139_p2 = (a0_389_fu_7756_p2 ^ a0_381_fu_7875_p2);

assign a0_386_fu_8155_p2 = (a0_390_fu_8129_p1 ^ a0_382_fu_7893_p2);

assign a0_387_fu_8235_p2 = (a0_388_fu_8221_p3 ^ a0_386_fu_8155_p2);

assign a0_388_fu_8221_p3 = a_259_fu_8133_p2[32'd2];

assign a0_389_fu_7756_p2 = (z2_192_fu_7716_p3 ^ z0_61_fu_7614_p3);

assign a0_390_fu_8129_p1 = a0_389_fu_7756_p2[0:0];

assign a0_391_fu_8461_p2 = (a0_392_fu_8451_p1 ^ a0_390_fu_8129_p1);

assign a0_392_fu_8451_p1 = a1_360_fu_7750_p2[0:0];

assign a0_393_fu_9245_p3 = {{a1_367_fu_9215_p2}, {a0_394_fu_9191_p2}};

assign a0_394_fu_9191_p2 = (z2_201_fu_9143_p3 ^ z0_85_fu_8841_p3);

assign a0_395_fu_9203_p2 = (xor_ln45_219_fu_8835_p2 ^ a0_206_fu_9137_p2);

assign a0_396_fu_9233_p2 = (xor_ln43_fu_9221_p2 ^ xor_ln43_71_fu_9227_p2);

assign a0_397_fu_9354_p2 = (a0_398_fu_9340_p3 ^ a0_396_fu_9233_p2);

assign a0_398_fu_9340_p3 = a0_394_fu_9191_p2[32'd2];

assign a0_399_fu_9523_p2 = (a0_403_fu_9519_p1 ^ a0_395_fu_9203_p2);

assign a0_400_fu_9539_p2 = (a0_404_fu_9515_p1 ^ a0_396_fu_9233_p2);

assign a0_401_fu_9619_p2 = (a0_402_fu_9605_p3 ^ a0_400_fu_9539_p2);

assign a0_402_fu_9605_p3 = a_309_fu_9197_p2[32'd2];

assign a0_403_fu_9519_p1 = a1_367_fu_9215_p2[1:0];

assign a0_404_fu_9515_p1 = a1_367_fu_9215_p2[0:0];

assign a0_405_fu_9859_p2 = (a0_406_fu_9845_p3 ^ a0_404_fu_9515_p1);

assign a0_406_fu_9845_p3 = a1_367_fu_9215_p2[32'd2];

assign a0_407_fu_10124_p2 = (a0_420_fu_8692_p2 ^ a0_394_fu_9191_p2);

assign a0_408_fu_10140_p2 = (a0_421_fu_10096_p1 ^ a0_395_fu_9203_p2);

assign a0_409_fu_10156_p2 = (a0_422_fu_10092_p1 ^ a0_396_fu_9233_p2);

assign a0_410_fu_10236_p2 = (a0_411_fu_10222_p3 ^ a0_409_fu_10156_p2);

assign a0_411_fu_10222_p3 = a0_407_fu_10124_p2[32'd2];

assign a0_412_fu_10427_p2 = (a0_416_fu_10411_p4 ^ a0_408_fu_10140_p2);

assign a0_413_fu_10443_p2 = (a0_417_fu_10403_p3 ^ a0_409_fu_10156_p2);

assign a0_414_fu_10524_p2 = (a0_415_fu_10510_p3 ^ a0_413_fu_10443_p2);

assign a0_415_fu_10510_p3 = a_354_fu_10421_p2[32'd2];

assign a0_416_fu_10411_p4 = {{a_339_fu_10112_p2[5:4]}};

assign a0_417_fu_10403_p3 = a_339_fu_10112_p2[32'd4];

assign a0_418_fu_10769_p2 = (a0_419_fu_10755_p3 ^ a0_417_fu_10403_p3);

assign a0_419_cast_fu_9253_p3 = {{xor_ln45_306_fu_9239_p2}, {a0_394_fu_9191_p2}};

assign a0_419_fu_10755_p3 = a_339_fu_10112_p2[32'd6];

assign a0_420_fu_8692_p2 = (z2_197_fu_8614_p3 ^ z0_72_fu_8121_p3);

assign a0_421_fu_10096_p1 = a0_420_fu_8692_p2[1:0];

assign a0_422_fu_10092_p1 = a0_420_fu_8692_p2[0:0];

assign a0_423_fu_11080_p2 = (a0_424_fu_11066_p3 ^ a0_422_fu_10092_p1);

assign a0_424_fu_11066_p3 = a0_420_fu_8692_p2[32'd2];

assign a0_425_fu_11251_p2 = (a0_429_fu_10100_p1 ^ a0_421_fu_10096_p1);

assign a0_426_fu_11267_p2 = (a0_430_fu_11241_p1 ^ a0_422_fu_10092_p1);

assign a0_427_fu_11347_p2 = (a0_428_fu_11333_p3 ^ a0_426_fu_11267_p2);

assign a0_428_fu_11333_p3 = a_399_fu_11245_p2[32'd2];

assign a0_429_fu_10100_p1 = a1_395_fu_8686_p2[1:0];

assign a0_430_fu_11241_p1 = a1_395_fu_8686_p2[0:0];

assign a0_431_fu_11587_p2 = (a0_432_fu_11573_p3 ^ a0_430_fu_11241_p1);

assign a0_432_fu_11573_p3 = a1_395_fu_8686_p2[32'd2];

assign a0_45_fu_2400_p2 = (z2_19_fu_2388_p2 ^ z0_22_fu_2364_p2);

assign a0_49_fu_2704_p2 = (z2_23_fu_2692_p2 ^ z0_26_fu_2668_p2);

assign a0_50_fu_2750_p2 = (z2_180_fu_2710_p3 ^ z0_24_fu_2538_p3);

assign a0_52_fu_2764_p1 = a1_290_fu_2744_p2[0:0];

assign a0_57_fu_3124_p2 = (z2_28_fu_3112_p2 ^ z0_30_fu_3088_p2);

assign a0_64_fu_3500_p2 = (z2_32_fu_3488_p2 ^ z0_35_fu_3464_p2);

assign a0_69_fu_3804_p2 = (z2_36_fu_3792_p2 ^ z0_39_fu_3768_p2);

assign a0_70_fu_3850_p2 = (z2_184_fu_3810_p3 ^ z0_37_fu_3638_p3);

assign a0_72_fu_3864_p1 = a1_304_fu_3844_p2[0:0];

assign a0_73_fu_3934_p2 = (z2_185_fu_3856_p3 ^ z0_31_fu_3176_p3);

assign a0_74_fu_3960_p1 = a1_305_fu_3928_p2[1:0];

assign a0_76_fu_3974_p3 = a1_305_fu_3928_p2[32'd2];

assign a0_86_fu_4300_p2 = (a1_sqr_25_fu_4292_p3 ^ a0_sqr_5_fu_4262_p3);

assign a0_94_fu_4468_p2 = (a1_sqr_28_fu_4460_p3 ^ a0_sqr_13_fu_4452_p3);

assign a0_96_fu_4506_p2 = (a1_sqr_29_fu_4484_p3 ^ a0_sqr_11_fu_4422_p3);

assign a0_98_fu_4522_p1 = a1_315_fu_4500_p2[0:0];

assign a0_fu_788_p2 = (z2_2_fu_776_p2 ^ z0_3_fu_752_p2);

assign a0_sqr_11_fu_4422_p3 = {{tmp_217_fu_4412_p4}, {xor_ln59_9_fu_4406_p2}};

assign a0_sqr_13_fu_4452_p3 = {{a1_313_fu_4438_p3}, {b_344_fu_4446_p2}};

assign a0_sqr_16_fu_6628_p3 = {{a1_333_reg_14371}, {b_198_fu_6624_p2}};

assign a0_sqr_18_fu_6652_p3 = {{tmp_256_reg_14392}, {xor_ln59_16_fu_6646_p2}};

assign a0_sqr_1_fu_4178_p3 = {{a1_307_fu_4164_p3}, {b_238_fu_4172_p2}};

assign a0_sqr_20_fu_6663_p3 = {{a1_335_reg_14397}, {b_224_fu_6659_p2}};

assign a0_sqr_23_fu_7228_p3 = {{a1_342_fu_7214_p3}, {b_185_fu_7222_p2}};

assign a0_sqr_3_fu_4232_p3 = {{tmp_208_fu_4222_p4}, {xor_ln59_2_fu_4216_p2}};

assign a0_sqr_5_fu_4262_p3 = {{a1_309_fu_4248_p3}, {b_264_fu_4256_p2}};

assign a0_sqr_7_fu_4344_p4 = {{{xor_ln28_25_fu_4332_p2}, {tmp_213_fu_4306_p4}}, {xor_ln59_6_fu_4338_p2}};

assign a0_sqr_9_fu_4368_p3 = {{a1_311_fu_4354_p3}, {b_318_fu_4362_p2}};

assign a0z1_1_fu_4978_p2 = (tmp_29_fu_4830_p3 ^ a0_340_fu_4704_p2);

assign a0z1_2_fu_6872_p2 = (tmp_39_fu_6805_p3 ^ a0_362_fu_6743_p2);

assign a0z1_3_fu_7350_p2 = (tmp_43_fu_7342_p3 ^ a0_371_fu_7314_p2);

assign a0z1_4_fu_7456_p2 = (a1_345_fu_7448_p3 ^ a0_374_fu_7442_p2);

assign a0z1_fu_440_p2 = (tmp_3_fu_388_p3 ^ a0_284_fu_168_p1);

assign a1_103_fu_6284_p2 = (z1_47_fu_6274_p2 ^ z0_48_fu_6262_p2);

assign a1_109_fu_6468_p2 = (z1_52_fu_6458_p2 ^ z0_52_fu_6446_p2);

assign a1_111_fu_6538_p3 = a1_332_fu_6514_p2[32'd1];

assign a1_126_fu_7128_p2 = (z1_56_fu_7116_p2 ^ z0_56_fu_7098_p2);

assign a1_13_fu_782_p2 = (z1_3_fu_770_p2 ^ z0_3_fu_752_p2);

assign a1_141_fu_7704_p2 = (z1_63_fu_7696_p2 ^ z0_63_fu_7692_p2);

assign a1_142_fu_7841_p2 = (z1_67_fu_7833_p2 ^ z0_67_fu_7829_p2);

assign a1_149_fu_8063_p2 = (z1_71_fu_8053_p2 ^ z0_71_fu_8042_p2);

assign a1_155_fu_8336_p2 = (z1_75_fu_8325_p2 ^ z0_76_fu_8310_p2);

assign a1_161_fu_8556_p2 = (z1_80_fu_8546_p2 ^ z0_80_fu_8535_p2);

assign a1_163_fu_8626_p3 = a1_364_fu_8602_p2[32'd1];

assign a1_164_fu_8783_p2 = (z1_84_fu_8773_p2 ^ z0_84_fu_8768_p2);

assign a1_165_fu_8934_p2 = (z1_88_fu_8924_p2 ^ z0_89_fu_8919_p2);

assign a1_167_fu_9085_p2 = (z1_93_fu_9075_p2 ^ z0_93_fu_9070_p2);

assign a1_169_fu_9155_p3 = a1_365_fu_9131_p2[32'd1];

assign a1_178_fu_9449_p2 = (z1_97_fu_9439_p2 ^ z0_97_fu_9428_p2);

assign a1_183_fu_9720_p2 = (z1_101_fu_9709_p2 ^ z0_102_fu_9694_p2);

assign a1_190_fu_9954_p2 = (z1_106_fu_9944_p2 ^ z0_106_fu_9933_p2);

assign a1_192_fu_10024_p3 = a1_380_fu_10000_p2[32'd1];

assign a1_198_fu_10337_p2 = (z1_110_fu_10326_p2 ^ z0_111_fu_10311_p2);

assign a1_19_fu_1158_p2 = (z1_7_fu_1146_p2 ^ z0_8_fu_1128_p2);

assign a1_212_fu_10625_p2 = (z1_114_fu_10614_p2 ^ z0_116_fu_10599_p2);

assign a1_217_fu_10869_p2 = (z1_119_fu_10858_p2 ^ z0_120_fu_10843_p2);

assign a1_219_fu_10939_p3 = a1_394_fu_10915_p2[32'd1];

assign a1_225_fu_11175_p2 = (z1_124_fu_11165_p2 ^ z0_124_fu_11154_p2);

assign a1_230_fu_11448_p2 = (z1_128_fu_11437_p2 ^ z0_129_fu_11422_p2);

assign a1_236_fu_11752_p3 = a1_408_fu_11728_p2[32'd1];

assign a1_239_fu_11842_p3 = a1_409_fu_11800_p2[32'd3];

assign a1_240_fu_12001_p2 = (z1_137_fu_11991_p2 ^ z0_137_fu_11986_p2);

assign a1_241_fu_12152_p2 = (z1_141_fu_12142_p2 ^ z0_142_fu_12137_p2);

assign a1_242_fu_12303_p2 = (z1_146_fu_12293_p2 ^ z0_146_fu_12288_p2);

assign a1_244_fu_12373_p3 = a1_411_fu_12349_p2[32'd1];

assign a1_245_fu_12526_p2 = (z1_150_fu_12516_p2 ^ z0_151_fu_12511_p2);

assign a1_246_fu_12677_p2 = (z1_154_fu_12667_p2 ^ z0_156_fu_12662_p2);

assign a1_247_fu_12828_p2 = (z1_159_fu_12818_p2 ^ z0_160_fu_12813_p2);

assign a1_249_fu_12898_p3 = a1_412_fu_12874_p2[32'd1];

assign a1_24_fu_1462_p2 = (z1_12_fu_1450_p2 ^ z0_12_fu_1432_p2);

assign a1_250_fu_13051_p2 = (z1_164_fu_13041_p2 ^ z0_164_fu_13036_p2);

assign a1_251_fu_13202_p2 = (z1_168_fu_13192_p2 ^ z0_169_fu_13187_p2);

assign a1_252_fu_13353_p2 = (z1_173_fu_13343_p2 ^ z0_173_fu_13338_p2);

assign a1_254_fu_13423_p3 = a1_413_fu_13399_p2[32'd1];

assign a1_257_fu_13513_p3 = a1_414_fu_13471_p2[32'd3];

assign a1_258_fu_194_p4 = {{a[31:24]}};

assign a1_259_fu_214_p4 = {{a[31:28]}};

assign a1_260_fu_234_p4 = {{a[31:30]}};

assign a1_261_fu_252_p3 = a[32'd31];

assign a1_262_fu_464_p4 = {{a[15:8]}};

assign a1_263_fu_506_p4 = {{a[7:4]}};

assign a1_264_fu_532_p4 = {{a[3:2]}};

assign a1_265_fu_558_p3 = a[32'd1];

assign a1_266_fu_664_p3 = a_11_fu_638_p2[32'd1];

assign a1_267_fu_736_p3 = a[32'd3];

assign a1_268_fu_902_p4 = {{a_20_fu_866_p2[3:2]}};

assign a1_269_fu_934_p3 = a0_295_fu_896_p2[32'd1];

assign a1_270_fu_1040_p3 = a_25_fu_1014_p2[32'd1];

assign a1_271_fu_1112_p3 = a_20_fu_866_p2[32'd3];

assign a1_272_fu_1224_p4 = {{a[7:6]}};

assign a1_273_fu_1244_p3 = a[32'd5];

assign a1_274_fu_1344_p3 = a_39_fu_1318_p2[32'd1];

assign a1_275_fu_1416_p3 = a[32'd7];

assign a1_276_fu_1508_p2 = (xor_ln45_27_fu_1502_p2 ^ xor_ln45_26_fu_1496_p2);

assign a1_277_fu_1730_p4 = {{a_50_fu_1662_p2[7:4]}};

assign a1_278_fu_1762_p4 = {{a0_303_fu_1724_p2[3:2]}};

assign a1_279_fu_1794_p3 = a0_304_fu_1756_p2[32'd1];

assign a1_27_fu_1532_p3 = a1_276_fu_1508_p2[32'd1];

assign a1_280_fu_1900_p3 = a_56_fu_1874_p2[32'd1];

assign a1_281_fu_1972_p3 = a0_303_fu_1724_p2[32'd3];

assign a1_282_fu_2138_p4 = {{a_65_fu_2102_p2[3:2]}};

assign a1_283_fu_2170_p3 = a0_308_fu_2132_p2[32'd1];

assign a1_284_fu_2276_p3 = a_70_fu_2250_p2[32'd1];

assign a1_285_fu_2348_p3 = a_65_fu_2102_p2[32'd3];

assign a1_286_fu_2460_p4 = {{a_50_fu_1662_p2[7:6]}};

assign a1_287_fu_2480_p3 = xor_ln43_14_fu_1668_p2[32'd5];

assign a1_288_fu_2580_p3 = a_84_fu_2554_p2[32'd1];

assign a1_289_fu_2652_p3 = a_50_fu_1662_p2[32'd7];

assign a1_290_fu_2744_p2 = (xor_ln45_65_fu_2738_p2 ^ xor_ln45_64_fu_2732_p2);

assign a1_291_fu_2860_p4 = {{a[15:12]}};

assign a1_292_fu_2880_p4 = {{a[11:10]}};

assign a1_293_fu_2900_p3 = a[32'd9];

assign a1_294_fu_3000_p3 = a_101_fu_2974_p2[32'd1];

assign a1_295_fu_3072_p3 = a[32'd11];

assign a1_296_fu_3238_p4 = {{a_110_fu_3202_p2[3:2]}};

assign a1_297_fu_3270_p3 = a0_321_fu_3232_p2[32'd1];

assign a1_298_fu_3376_p3 = a_115_fu_3350_p2[32'd1];

assign a1_299_fu_3448_p3 = a_110_fu_3202_p2[32'd3];

assign a1_300_fu_3560_p4 = {{a[15:14]}};

assign a1_301_fu_3580_p3 = a[32'd13];

assign a1_302_fu_3680_p3 = a_129_fu_3654_p2[32'd1];

assign a1_303_fu_3752_p3 = a[32'd15];

assign a1_304_fu_3844_p2 = (xor_ln45_103_fu_3838_p2 ^ xor_ln45_102_fu_3832_p2);

assign a1_305_fu_3928_p2 = (xor_ln45_113_fu_3910_p2 ^ xor_ln45_112_fu_3904_p2);

assign a1_306_fu_3964_p4 = {{a1_305_fu_3928_p2[3:2]}};

assign a1_307_fu_4164_p3 = a[32'd17];

assign a1_308_fu_4194_p3 = a[32'd19];

assign a1_309_fu_4248_p3 = a[32'd21];

assign a1_310_fu_4278_p3 = a[32'd23];

assign a1_311_fu_4354_p3 = a[32'd25];

assign a1_312_fu_4384_p3 = a[32'd27];

assign a1_313_fu_4438_p3 = a[32'd29];

integer ap_tvar_int_0;

always @ (a) begin
    for (ap_tvar_int_0 = 2 - 1; ap_tvar_int_0 >= 0; ap_tvar_int_0 = ap_tvar_int_0 - 1) begin
        if (ap_tvar_int_0 > 31 - 30) begin
            a1_314_fu_4474_p4[ap_tvar_int_0] = 1'b0;
        end else begin
            a1_314_fu_4474_p4[ap_tvar_int_0] = a[31 - ap_tvar_int_0];
        end
    end
end

assign a1_315_fu_4500_p2 = (tmp_23_fu_4492_p3 ^ a0_94_fu_4468_p2);

assign a1_316_fu_4726_p4 = {{delta_fu_4668_p2[15:12]}};

assign a1_317_fu_4746_p4 = {{delta_fu_4668_p2[15:14]}};

assign a1_318_fu_4764_p3 = delta_fu_4668_p2[32'd15];

assign a1_319_fu_4990_p4 = {{a0_340_fu_4704_p2[7:4]}};

assign a1_320_fu_5016_p4 = {{a0_344_fu_4964_p2[3:2]}};

assign a1_324_fu_5178_p4 = {{a_170_fu_5142_p2[3:2]}};

assign a1_328_fu_5280_p4 = {{a0_340_fu_4704_p2[7:6]}};

assign a1_332_fu_6514_p2 = (xor_ln45_172_fu_6508_p2 ^ xor_ln45_171_fu_6502_p2);

assign a1_336_fu_6759_p4 = {{delta_1_fu_6731_p2[7:6]}};

assign a1_337_fu_6777_p3 = delta_1_fu_6731_p2[32'd7];

assign a1_338_fu_6878_p4 = {{a0_362_fu_6743_p2[3:2]}};

assign a1_339_fu_6904_p3 = a0_365_fu_6866_p2[32'd1];

assign a1_340_fu_7010_p3 = a_210_fu_6984_p2[32'd1];

assign a1_341_fu_7082_p3 = a0_362_fu_6743_p2[32'd3];

assign a1_342_fu_7214_p3 = xor_ln71_4_fu_6737_p2[32'd5];

assign a1_343_fu_7328_p3 = delta_2_fu_7284_p2[32'd3];

assign a1_344_fu_7362_p3 = a0_371_fu_7314_p2[32'd1];

assign a1_345_fu_7448_p3 = delta_3_fu_7436_p2[32'd1];

assign a1_346_fu_7474_p2 = (delta_4_fu_7468_p2 & a1_345_fu_7448_p3);

assign a1_347_fu_7584_p3 = {{a1_350_reg_14762}, {a0_379_reg_14769}};

assign a1_348_fu_7540_p2 = (z1_59_fu_7528_p2 ^ z0_59_fu_7522_p2);

assign a1_349_fu_7632_p3 = a_235_fu_7622_p2[32'd1];

assign a1_34_fu_2018_p2 = (z1_16_fu_2006_p2 ^ z0_17_fu_1988_p2);

assign a1_350_fu_7510_p2 = (z1_58_fu_7498_p2 ^ z0_58_fu_7486_p2);

assign a1_351_fu_7907_p3 = {{a1_360_fu_7750_p2}, {a0_389_fu_7756_p2}};

assign a1_352_fu_7887_p2 = (a_250_fu_7881_p2 ^ a0_381_fu_7875_p2);

assign a1_353_fu_7915_p3 = a0_381_fu_7875_p2[32'd1];

assign a1_354_fu_7974_p3 = a_250_fu_7881_p2[32'd1];

assign a1_355_fu_8034_p3 = a1_352_fu_7887_p2[32'd1];

assign a1_356_fu_8145_p4 = {{a_259_fu_8133_p2[3:2]}};

assign a1_357_fu_8161_p3 = a0_385_fu_8139_p2[32'd1];

assign a1_358_fu_8241_p3 = a_264_fu_8229_p2[32'd1];

assign a1_359_fu_8302_p3 = a_259_fu_8133_p2[32'd3];

assign a1_360_fu_7750_p2 = (xor_ln45_209_fu_7744_p2 ^ xor_ln45_208_fu_7738_p2);

assign a1_361_fu_8402_p3 = a0_389_fu_7756_p2[32'd1];

assign a1_362_fu_8467_p3 = a_278_fu_8455_p2[32'd1];

assign a1_363_fu_8527_p3 = a1_360_fu_7750_p2[32'd1];

assign a1_364_fu_8602_p2 = (xor_ln45_248_fu_8596_p2 ^ xor_ln45_243_fu_8590_p2);

assign a1_365_fu_9131_p2 = (xor_ln45_292_fu_9125_p2 ^ xor_ln45_285_fu_9119_p2);

assign a1_366_fu_9273_p3 = {{a1_395_fu_8686_p2}, {a0_420_fu_8692_p2}};

assign a1_367_fu_9215_p2 = (a_309_fu_9197_p2 ^ a0_394_fu_9191_p2);

assign a1_368_fu_9281_p4 = {{a0_394_fu_9191_p2[3:2]}};

assign a1_369_fu_9291_p3 = a0_395_fu_9203_p2[32'd1];

assign a1_370_fu_9360_p3 = a_300_fu_9348_p2[32'd1];

assign a1_371_fu_9420_p3 = a0_394_fu_9191_p2[32'd3];

assign a1_372_fu_9529_p4 = {{a_309_fu_9197_p2[3:2]}};

assign a1_373_fu_9545_p3 = a0_399_fu_9523_p2[32'd1];

assign a1_374_fu_9625_p3 = a_314_fu_9613_p2[32'd1];

assign a1_375_fu_9686_p3 = a_309_fu_9197_p2[32'd3];

assign a1_376_fu_9786_p4 = {{a1_367_fu_9215_p2[3:2]}};

assign a1_377_fu_9796_p3 = xor_ln45_306_fu_9239_p2[32'd1];

assign a1_378_fu_9865_p3 = a_328_fu_9853_p2[32'd1];

assign a1_379_fu_9925_p3 = a1_367_fu_9215_p2[32'd3];

assign a1_380_fu_10000_p2 = (xor_ln45_336_fu_9994_p2 ^ xor_ln45_329_fu_9988_p2);

assign a1_381_fu_10130_p4 = {{a_339_fu_10112_p2[7:4]}};

assign a1_382_fu_10146_p4 = {{a0_407_fu_10124_p2[3:2]}};

assign a1_383_fu_10162_p3 = a0_408_fu_10140_p2[32'd1];

assign a1_384_fu_10242_p3 = a_345_fu_10230_p2[32'd1];

assign a1_385_fu_10303_p3 = a0_407_fu_10124_p2[32'd3];

assign a1_386_fu_10433_p4 = {{a_354_fu_10421_p2[3:2]}};

assign a1_387_fu_10449_p3 = a0_412_fu_10427_p2[32'd1];

assign a1_388_fu_10530_p3 = a_359_fu_10518_p2[32'd1];

assign a1_389_fu_10591_p3 = a_354_fu_10421_p2[32'd3];

assign a1_390_fu_10691_p4 = {{a_339_fu_10112_p2[7:6]}};

assign a1_391_fu_10701_p3 = xor_ln43_83_fu_10118_p2[32'd5];

assign a1_392_fu_10775_p3 = a_373_fu_10763_p2[32'd1];

assign a1_393_fu_10835_p3 = a_339_fu_10112_p2[32'd7];

assign a1_394_fu_10915_p2 = (xor_ln45_364_fu_10909_p2 ^ xor_ln45_357_fu_10903_p2);

assign a1_395_fu_8686_p2 = (xor_ln45_258_fu_8668_p2 ^ xor_ln45_251_fu_8662_p2);

assign a1_396_fu_11007_p4 = {{a0_420_fu_8692_p2[3:2]}};

assign a1_397_fu_11017_p3 = xor_ln73_fu_9261_p2[32'd1];

assign a1_398_fu_11086_p3 = a_390_fu_11074_p2[32'd1];

assign a1_399_fu_11146_p3 = a0_420_fu_8692_p2[32'd3];

assign a1_400_fu_11257_p4 = {{a_399_fu_11245_p2[3:2]}};

assign a1_401_fu_11273_p3 = a0_425_fu_11251_p2[32'd1];

assign a1_402_fu_11353_p3 = a_404_fu_11341_p2[32'd1];

assign a1_403_fu_11414_p3 = a_399_fu_11245_p2[32'd3];

assign a1_404_fu_11514_p4 = {{a1_395_fu_8686_p2[3:2]}};

assign a1_405_fu_11524_p3 = xor_ln73_1_fu_9267_p2[32'd1];

assign a1_406_fu_11593_p3 = a_418_fu_11581_p2[32'd1];

assign a1_407_fu_11653_p3 = a1_395_fu_8686_p2[32'd3];

assign a1_408_fu_11728_p2 = (xor_ln45_398_fu_11722_p2 ^ xor_ln45_391_fu_11716_p2);

assign a1_409_fu_11800_p2 = (xor_ln45_408_fu_11794_p2 ^ xor_ln45_401_fu_11788_p2);

assign a1_40_fu_2394_p2 = (z1_20_fu_2382_p2 ^ z0_22_fu_2364_p2);

assign a1_410_fu_11824_p4 = {{a1_409_fu_11800_p2[3:2]}};

assign a1_411_fu_12349_p2 = (xor_ln45_442_fu_12343_p2 ^ xor_ln45_435_fu_12337_p2);

assign a1_412_fu_12874_p2 = (xor_ln45_460_fu_12868_p2 ^ xor_ln45_459_fu_12862_p2);

assign a1_413_fu_13399_p2 = (xor_ln45_476_fu_13393_p2 ^ xor_ln45_475_fu_13387_p2);

assign a1_414_fu_13471_p2 = (xor_ln45_480_fu_13465_p2 ^ xor_ln45_479_fu_13459_p2);

assign a1_415_fu_13495_p4 = {{a1_414_fu_13471_p2[3:2]}};

assign a1_46_fu_2698_p2 = (z1_25_fu_2686_p2 ^ z0_26_fu_2668_p2);

assign a1_49_fu_2768_p3 = a1_290_fu_2744_p2[32'd1];

assign a1_56_fu_3118_p2 = (z1_30_fu_3106_p2 ^ z0_30_fu_3088_p2);

assign a1_61_fu_3494_p2 = (z1_34_fu_3482_p2 ^ z0_35_fu_3464_p2);

assign a1_66_fu_3798_p2 = (z1_39_fu_3786_p2 ^ z0_39_fu_3768_p2);

assign a1_68_fu_3868_p3 = a1_304_fu_3844_p2[32'd1];

assign a1_71_fu_3982_p3 = a1_305_fu_3928_p2[32'd3];

assign a1_88_fu_4526_p3 = a1_315_fu_4500_p2[32'd1];

assign a1_98_fu_6086_p2 = (z1_43_fu_6076_p2 ^ z0_43_fu_6064_p2);

assign a1_fu_11682_p2 = (z1_133_fu_11672_p2 ^ z0_133_fu_11661_p2);

assign a1_sqr_25_fu_4292_p3 = {{a1_310_fu_4278_p3}, {a0_334_fu_4286_p2}};

assign a1_sqr_26_fu_4316_p3 = {{tmp_213_fu_4306_p4}, {a0_86_fu_4300_p2}};

assign a1_sqr_27_fu_4398_p3 = {{a1_312_fu_4384_p3}, {a0_337_fu_4392_p2}};

assign a1_sqr_28_fu_4460_p3 = {{a1_261_fu_252_p3}, {a0_339_fu_260_p2}};

assign a1_sqr_29_fu_4484_p3 = {{a1_314_fu_4474_p4}, {a0_94_fu_4468_p2}};

assign a1_sqr_30_fu_4512_p4 = {{{a1_315_fu_4500_p2}, {a1_314_fu_4474_p4}}, {a0_96_fu_4506_p2}};

assign a1_sqr_31_fu_6639_p3 = {{a1_334_reg_14385}, {a0_359_fu_6635_p2}};

assign a1_sqr_32_fu_6670_p3 = {{a1_318_reg_14145}, {a0_361_reg_14151}};

assign a1_sqr_33_fu_6682_p3 = {{tmp_258_reg_14404}, {a0_138_fu_6676_p2}};

assign a1_sqr_34_fu_7236_p3 = {{a1_337_fu_6777_p3}, {a0_370_fu_6785_p2}};

assign a1_sqr_fu_4208_p3 = {{a1_308_fu_4194_p3}, {a0_331_fu_4202_p2}};

assign a_101_fu_2974_p2 = (a1_292_fu_2880_p4 ^ a0_317_fu_1632_p4);

assign a_103_fu_3028_p2 = (a1_294_fu_3000_p3 ^ a0_319_fu_2994_p2);

assign a_107_fu_3094_p2 = (a1_295_fu_3072_p3 ^ a0_320_fu_2966_p3);

assign a_110_fu_3202_p2 = (a1_291_fu_2860_p4 ^ a0_316_fu_1642_p4);

assign a_113_fu_3298_p2 = (a1_297_fu_3270_p3 ^ a0_322_fu_3264_p2);

assign a_115_fu_3350_p2 = (a1_296_fu_3238_p4 ^ a0_321_fu_3232_p2);

assign a_117_fu_3404_p2 = (a1_298_fu_3376_p3 ^ a0_323_fu_3370_p2);

assign a_11_fu_638_p2 = (a1_264_fu_532_p4 ^ a0_291_fu_400_p1);

assign a_121_fu_3470_p2 = (a1_299_fu_3448_p3 ^ a0_324_fu_3342_p3);

assign a_127_fu_3602_p2 = (a1_301_fu_3580_p3 ^ a0_326_fu_3184_p3);

assign a_129_fu_3654_p2 = (a1_300_fu_3560_p4 ^ a0_325_fu_3192_p4);

assign a_131_fu_3708_p2 = (a1_302_fu_3680_p3 ^ a0_327_fu_3674_p2);

assign a_135_fu_3774_p2 = (a1_303_fu_3752_p3 ^ a0_328_fu_3646_p3);

assign a_13_fu_692_p2 = (a1_266_fu_664_p3 ^ a0_293_fu_658_p2);

assign a_159_fu_5972_p2 = (a1_321_reg_14175 ^ a0_346_reg_14167);

assign a_161_fu_5072_p2 = (a1_320_fu_5016_p4 ^ a0_345_fu_4946_p2);

assign a_163_fu_6024_p2 = (a1_322_reg_14212 ^ a0_347_fu_6010_p2);

assign a_167_fu_6068_p2 = (a1_323_reg_14225 ^ a0_348_reg_14197);

assign a_170_fu_5142_p2 = (a1_319_fu_4990_p4 ^ a0_344_fu_4964_p2);

assign a_173_fu_6166_p2 = (a1_325_reg_14255 ^ a0_350_fu_6152_p2);

assign a_175_fu_5228_p2 = (a1_324_fu_5178_p4 ^ a0_349_fu_5172_p2);

assign a_177_fu_6222_p2 = (a1_326_reg_14283 ^ a0_351_fu_6206_p2);

assign a_17_fu_758_p2 = (a1_267_fu_736_p3 ^ a0_294_fu_630_p3);

assign a_181_fu_6266_p2 = (a1_327_reg_14296 ^ a0_352_reg_14268);

assign a_187_fu_6354_p2 = (a1_329_reg_14309 ^ a0_354_reg_14238);

assign a_189_fu_5324_p2 = (a1_328_fu_5280_p4 ^ a0_353_fu_5132_p4);

assign a_191_fu_6406_p2 = (a1_330_reg_14337 ^ a0_355_fu_6392_p2);

assign a_195_fu_6450_p2 = (a1_331_reg_14350 ^ a0_356_reg_14322);

assign a_208_fu_6932_p2 = (a1_339_fu_6904_p3 ^ a0_366_fu_6848_p2);

assign a_20_fu_866_p2 = (a1_263_fu_506_p4 ^ a0_290_fu_404_p1);

assign a_210_fu_6984_p2 = (a1_338_fu_6878_p4 ^ a0_365_fu_6866_p2);

assign a_212_fu_7038_p2 = (a1_340_fu_7010_p3 ^ a0_367_fu_7004_p2);

assign a_216_fu_7104_p2 = (a1_341_fu_7082_p3 ^ a0_368_fu_6976_p3);

assign a_223_fu_7384_p2 = (a1_344_fu_7362_p3 ^ a0_373_fu_7308_p2);

assign a_229_fu_7492_p2 = (delta_4_fu_7468_p2 & a0_374_fu_7442_p2);

assign a_233_fu_7552_p2 = (z2_59_fu_7534_p2 ^ z1_59_fu_7528_p2);

assign a_235_fu_7622_p2 = (a1_347_fu_7584_p3 ^ a0_376_fu_7578_p3);

assign a_237_fu_7650_p2 = (a1_349_fu_7632_p3 ^ a0_378_fu_7628_p2);

assign a_23_fu_962_p2 = (a1_269_fu_934_p3 ^ a0_296_fu_928_p2);

assign a_241_fu_7572_p2 = (z2_58_fu_7504_p2 ^ z1_58_fu_7498_p2);

assign a_248_fu_7928_p2 = (a1_353_fu_7915_p3 ^ a0_382_fu_7893_p2);

assign a_250_fu_7881_p2 = (z1_66_fu_7821_p3 ^ tmp_47_fu_7867_p3);

assign a_252_fu_7992_p2 = (a1_354_fu_7974_p3 ^ a0_383_fu_7968_p2);

assign a_256_fu_8047_p2 = (a1_355_fu_8034_p3 ^ a0_384_fu_7964_p1);

assign a_259_fu_8133_p2 = (a1_351_fu_7907_p3 ^ a0_380_fu_7899_p3);

assign a_25_fu_1014_p2 = (a1_268_fu_902_p4 ^ a0_295_fu_896_p2);

assign a_262_fu_8179_p2 = (a1_357_fu_8161_p3 ^ a0_386_fu_8155_p2);

assign a_264_fu_8229_p2 = (a1_356_fu_8145_p4 ^ a0_385_fu_8139_p2);

assign a_266_fu_8260_p2 = (a1_358_fu_8241_p3 ^ a0_387_fu_8235_p2);

assign a_270_fu_8315_p2 = (a1_359_fu_8302_p3 ^ a0_388_fu_8221_p3);

assign a_276_fu_8415_p2 = (a1_361_fu_8402_p3 ^ a0_390_fu_8129_p1);

assign a_278_fu_8455_p2 = (a1_360_fu_7750_p2 ^ a0_389_fu_7756_p2);

assign a_27_fu_1068_p2 = (a1_270_fu_1040_p3 ^ a0_297_fu_1034_p2);

assign a_280_fu_8485_p2 = (a1_362_fu_8467_p3 ^ a0_391_fu_8461_p2);

assign a_284_fu_8540_p2 = (a1_363_fu_8527_p3 ^ a0_392_fu_8451_p1);

assign a_298_fu_9304_p2 = (a1_369_fu_9291_p3 ^ a0_396_fu_9233_p2);

assign a_300_fu_9348_p2 = (a1_368_fu_9281_p4 ^ a0_395_fu_9203_p2);

assign a_302_fu_9378_p2 = (a1_370_fu_9360_p3 ^ a0_397_fu_9354_p2);

assign a_306_fu_9433_p2 = (a1_371_fu_9420_p3 ^ a0_398_fu_9340_p3);

assign a_309_fu_9197_p2 = (z1_89_fu_8992_p3 ^ tmp_57_fu_9183_p3);

assign a_312_fu_9563_p2 = (a1_373_fu_9545_p3 ^ a0_400_fu_9539_p2);

assign a_314_fu_9613_p2 = (a1_372_fu_9529_p4 ^ a0_399_fu_9523_p2);

assign a_316_fu_9644_p2 = (a1_374_fu_9625_p3 ^ a0_401_fu_9619_p2);

assign a_31_fu_1134_p2 = (a1_271_fu_1112_p3 ^ a0_298_fu_1006_p3);

assign a_320_fu_9699_p2 = (a1_375_fu_9686_p3 ^ a0_402_fu_9605_p3);

assign a_326_fu_9809_p2 = (a1_377_fu_9796_p3 ^ a0_404_fu_9515_p1);

assign a_328_fu_9853_p2 = (a1_376_fu_9786_p4 ^ a0_403_fu_9519_p1);

assign a_330_fu_9883_p2 = (a1_378_fu_9865_p3 ^ a0_405_fu_9859_p2);

assign a_334_fu_9938_p2 = (a1_379_fu_9925_p3 ^ a0_406_fu_9845_p3);

assign a_339_fu_10112_p2 = (a1_366_fu_9273_p3 ^ a0_393_fu_9245_p3);

assign a_343_fu_10180_p2 = (a1_383_fu_10162_p3 ^ a0_409_fu_10156_p2);

assign a_345_fu_10230_p2 = (a1_382_fu_10146_p4 ^ a0_408_fu_10140_p2);

assign a_347_fu_10261_p2 = (a1_384_fu_10242_p3 ^ a0_410_fu_10236_p2);

assign a_351_fu_10316_p2 = (a1_385_fu_10303_p3 ^ a0_411_fu_10222_p3);

assign a_354_fu_10421_p2 = (a1_381_fu_10130_p4 ^ a0_407_fu_10124_p2);

assign a_357_fu_10468_p2 = (a1_387_fu_10449_p3 ^ a0_413_fu_10443_p2);

assign a_359_fu_10518_p2 = (a1_386_fu_10433_p4 ^ a0_412_fu_10427_p2);

assign a_361_fu_10549_p2 = (a1_388_fu_10530_p3 ^ a0_414_fu_10524_p2);

assign a_365_fu_10604_p2 = (a1_389_fu_10591_p3 ^ a0_415_fu_10510_p3);

assign a_371_fu_10714_p2 = (a1_391_fu_10701_p3 ^ a0_417_fu_10403_p3);

assign a_373_fu_10763_p2 = (a1_390_fu_10691_p4 ^ a0_416_fu_10411_p4);

assign a_375_fu_10793_p2 = (a1_392_fu_10775_p3 ^ a0_418_fu_10769_p2);

assign a_379_fu_10848_p2 = (a1_393_fu_10835_p3 ^ a0_419_fu_10755_p3);

assign a_37_fu_1266_p2 = (a1_273_fu_1244_p3 ^ a0_300_fu_848_p3);

assign a_388_fu_11030_p2 = (a1_397_fu_11017_p3 ^ a0_422_fu_10092_p1);

assign a_390_fu_11074_p2 = (a1_396_fu_11007_p4 ^ a0_421_fu_10096_p1);

assign a_392_fu_11104_p2 = (a1_398_fu_11086_p3 ^ a0_423_fu_11080_p2);

assign a_396_fu_11159_p2 = (a1_399_fu_11146_p3 ^ a0_424_fu_11066_p3);

assign a_399_fu_11245_p2 = (a1_395_fu_8686_p2 ^ a0_420_fu_8692_p2);

assign a_39_fu_1318_p2 = (a1_272_fu_1224_p4 ^ a0_299_fu_856_p4);

assign a_402_fu_11291_p2 = (a1_401_fu_11273_p3 ^ a0_426_fu_11267_p2);

assign a_404_fu_11341_p2 = (a1_400_fu_11257_p4 ^ a0_425_fu_11251_p2);

assign a_406_fu_11372_p2 = (a1_402_fu_11353_p3 ^ a0_427_fu_11347_p2);

assign a_410_fu_11427_p2 = (a1_403_fu_11414_p3 ^ a0_428_fu_11333_p3);

assign a_416_fu_11537_p2 = (a1_405_fu_11524_p3 ^ a0_430_fu_11241_p1);

assign a_418_fu_11581_p2 = (a1_404_fu_11514_p4 ^ a0_429_fu_10100_p1);

assign a_41_fu_1372_p2 = (a1_274_fu_1344_p3 ^ a0_301_fu_1338_p2);

assign a_420_fu_11611_p2 = (a1_406_fu_11593_p3 ^ a0_431_fu_11587_p2);

assign a_424_fu_11666_p2 = (a1_407_fu_11653_p3 ^ a0_432_fu_11573_p3);

assign a_45_fu_1438_p2 = (a1_275_fu_1416_p3 ^ a0_302_fu_1310_p3);

assign a_50_fu_1662_p2 = (a1_262_fu_464_p4 ^ a0_289_fu_408_p1);

assign a_54_fu_1822_p2 = (a1_279_fu_1794_p3 ^ a0_305_fu_1788_p2);

assign a_56_fu_1874_p2 = (a1_278_fu_1762_p4 ^ a0_304_fu_1756_p2);

assign a_58_fu_1928_p2 = (a1_280_fu_1900_p3 ^ a0_306_fu_1894_p2);

assign a_62_fu_1994_p2 = (a1_281_fu_1972_p3 ^ a0_307_fu_1866_p3);

assign a_65_fu_2102_p2 = (a1_277_fu_1730_p4 ^ a0_303_fu_1724_p2);

assign a_68_fu_2198_p2 = (a1_283_fu_2170_p3 ^ a0_309_fu_2164_p2);

assign a_70_fu_2250_p2 = (a1_282_fu_2138_p4 ^ a0_308_fu_2132_p2);

assign a_72_fu_2304_p2 = (a1_284_fu_2276_p3 ^ a0_310_fu_2270_p2);

assign a_76_fu_2370_p2 = (a1_285_fu_2348_p3 ^ a0_311_fu_2242_p3);

assign a_82_fu_2502_p2 = (a1_287_fu_2480_p3 ^ a0_313_fu_2084_p3);

assign a_84_fu_2554_p2 = (a1_286_fu_2460_p4 ^ a0_312_fu_2092_p4);

assign a_86_fu_2608_p2 = (a1_288_fu_2580_p3 ^ a0_314_fu_2574_p2);

assign a_90_fu_2674_p2 = (a1_289_fu_2652_p3 ^ a0_315_fu_2546_p3);

assign a_99_fu_2922_p2 = (a1_293_fu_2900_p3 ^ a0_318_fu_1624_p3);

assign a_9_fu_586_p2 = (a1_265_fu_558_p3 ^ a0_292_fu_396_p1);

assign and_ln36_fu_7462_p2 = (a0z1_4_fu_7456_p2 & a0_374_fu_7442_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_return = {{{{xor_ln45_348_fu_11904_p2}, {xor_ln45_349_fu_11910_p2}}, {xor_ln45_454_fu_13575_p2}}, {xor_ln45_455_fu_13581_p2}};

assign b0_10_fu_880_p4 = {{b0_fu_484_p2[5:4]}};

assign b0_11_fu_872_p3 = b0_fu_484_p2[32'd4];

assign b0_12_fu_1352_p2 = (b0_13_fu_1324_p3 ^ b0_11_fu_872_p3);

assign b0_13_fu_1324_p3 = b0_fu_484_p2[32'd6];

assign b0_14_fu_1740_p2 = (b0_27_fu_1692_p4 ^ b0_1_fu_516_p2);

assign b0_15_fu_1772_p2 = (b0_2_fu_542_p2 ^ b0_28_fu_1682_p4);

assign b0_16_fu_1802_p2 = (b0_3_fu_566_p2 ^ b0_29_fu_1674_p3);

assign b0_17_fu_1908_p2 = (b0_18_fu_1880_p3 ^ b0_16_fu_1802_p2);

assign b0_18_fu_1880_p3 = b0_14_fu_1740_p2[32'd2];

assign b0_19_fu_2148_p2 = (b0_23_fu_2116_p4 ^ b0_15_fu_1772_p2);

assign b0_1_fu_516_p2 = (a0_290_fu_404_p1 ^ a0_286_fu_204_p4);

assign b0_20_fu_2178_p2 = (b0_24_fu_2108_p3 ^ b0_16_fu_1802_p2);

assign b0_21_fu_2284_p2 = (b0_22_fu_2256_p3 ^ b0_20_fu_2178_p2);

assign b0_22_fu_2256_p3 = b_55_fu_2126_p2[32'd2];

assign b0_23_fu_2116_p4 = {{b_41_fu_1712_p2[5:4]}};

assign b0_24_fu_2108_p3 = b_41_fu_1712_p2[32'd4];

assign b0_25_fu_2588_p2 = (b0_26_fu_2560_p3 ^ b0_24_fu_2108_p3);

assign b0_26_fu_2560_p3 = b_41_fu_1712_p2[32'd6];

assign b0_27_fu_1692_p4 = {{a0z1_fu_440_p2[11:8]}};

assign b0_28_fu_1682_p4 = {{a0z1_fu_440_p2[9:8]}};

assign b0_29_fu_1674_p3 = a0z1_fu_440_p2[32'd8];

assign b0_2_fu_542_p2 = (b0_88_fu_288_p4 ^ a0_291_fu_400_p1);

assign b0_30_fu_3008_p2 = (b0_31_fu_2980_p3 ^ b0_29_fu_1674_p3);

assign b0_31_fu_2980_p3 = xor_ln70_3_fu_458_p2[32'd10];

assign b0_32_fu_3248_p2 = (b0_36_fu_3216_p4 ^ b0_28_fu_1682_p4);

assign b0_33_fu_3278_p2 = (b0_37_fu_3208_p3 ^ b0_29_fu_1674_p3);

assign b0_34_fu_3384_p2 = (b0_35_fu_3356_p3 ^ b0_33_fu_3278_p2);

assign b0_35_fu_3356_p3 = b_95_fu_3226_p2[32'd2];

assign b0_36_fu_3216_p4 = {{a0z1_fu_440_p2[13:12]}};

assign b0_37_fu_3208_p3 = a0z1_fu_440_p2[32'd12];

assign b0_38_fu_3688_p2 = (b0_39_fu_3660_p3 ^ b0_37_fu_3208_p3);

assign b0_39_fu_3660_p3 = a0z1_fu_440_p2[32'd14];

assign b0_3_fu_566_p2 = (a0_335_fu_362_p3 ^ a0_292_fu_396_p1);

assign b0_40_fu_5000_p2 = (a1_316_fu_4726_p4 ^ a0_344_fu_4964_p2);

assign b0_41_fu_5026_p2 = (a0_345_fu_4946_p2 ^ a0_342_fu_4736_p4);

assign b0_42_fu_5050_p2 = (a0_360_fu_4816_p3 ^ a0_346_fu_4922_p2);

assign b0_43_fu_6014_p2 = (b0_44_reg_14204 ^ b0_42_reg_14181);

assign b0_45_fu_5188_p2 = (b0_49_fu_5156_p4 ^ b0_41_fu_5026_p2);

assign b0_46_fu_6156_p2 = (b0_50_reg_14246 ^ b0_42_reg_14181);

assign b0_47_fu_6211_p2 = (b0_48_reg_14275 ^ b0_46_fu_6156_p2);

assign b0_49_fu_5156_p4 = {{a0z1_1_fu_4978_p2[5:4]}};

assign b0_4_fu_672_p2 = (b0_5_fu_644_p3 ^ b0_3_fu_566_p2);

assign b0_51_fu_6396_p2 = (b0_52_reg_14329 ^ b0_50_reg_14246);

assign b0_53_fu_6888_p2 = (a1_336_fu_6759_p4 ^ a0_365_fu_6866_p2);

assign b0_54_fu_6912_p2 = (a0_366_fu_6848_p2 ^ a0_364_fu_6769_p3);

assign b0_55_fu_7018_p2 = (b0_56_fu_6990_p3 ^ b0_54_fu_6912_p2);

assign b0_56_fu_6990_p3 = a0z1_2_fu_6872_p2[32'd2];

assign b0_57_fu_7356_p2 = (a1_343_fu_7328_p3 ^ a0_373_fu_7308_p2);

assign b0_58_fu_7640_p2 = (a0_369_reg_14746 ^ a0_364_reg_14685);

assign b0_59_fu_4800_p4 = {{xor_ln71_3_fu_4686_p2[9:8]}};

assign b0_5_fu_644_p3 = b0_1_fu_516_p2[32'd2];

assign b0_60_fu_7982_p2 = (a0_358_reg_14378_pp0_iter1_reg ^ a0_357_reg_14363_pp0_iter1_reg);

assign b0_61_fu_5466_p2 = (b0_59_fu_4800_p4 ^ a0_342_fu_4736_p4);

assign b0_62_fu_8169_p2 = (a0_360_reg_14159_pp0_iter1_reg ^ a0_357_reg_14363_pp0_iter1_reg);

assign b0_63_fu_8249_p2 = (b0_64_reg_14423_pp0_iter1_reg ^ b0_62_fu_8169_p2);

assign b0_65_fu_8475_p2 = (a0_360_reg_14159_pp0_iter1_reg ^ a0_343_reg_14138_pp0_iter1_reg);

assign b0_66_fu_318_p4 = {{a[19:16]}};

assign b0_67_fu_328_p4 = {{a[17:16]}};

assign b0_68_fu_9368_p2 = (a0_330_reg_14046_pp0_iter1_reg ^ a0_329_reg_14028_pp0_iter1_reg);

assign b0_69_fu_5584_p2 = (b0_73_fu_5568_p4 ^ b0_67_fu_328_p4);

assign b0_6_fu_912_p2 = (b0_2_fu_542_p2 ^ b0_10_fu_880_p4);

assign b0_70_fu_9553_p2 = (a0_332_reg_14062_pp0_iter1_reg ^ a0_329_reg_14028_pp0_iter1_reg);

assign b0_71_fu_9633_p2 = (b0_72_reg_14460_pp0_iter1_reg ^ b0_70_fu_9553_p2);

assign b0_73_fu_5568_p4 = {{a[21:20]}};

assign b0_74_fu_9873_p2 = (a0_333_reg_14079_pp0_iter1_reg ^ a0_332_reg_14062_pp0_iter1_reg);

assign b0_75_fu_5674_p2 = (b0_66_fu_318_p4 ^ a0_286_fu_204_p4);

assign b0_76_fu_5690_p2 = (b0_88_fu_288_p4 ^ b0_67_fu_328_p4);

assign b0_77_fu_10170_p2 = (a0_335_reg_13615_pp0_iter1_reg ^ a0_329_reg_14028_pp0_iter1_reg);

assign b0_78_fu_10250_p2 = (b0_79_reg_14491_pp0_iter1_reg ^ b0_77_fu_10170_p2);

assign b0_7_fu_942_p2 = (b0_3_fu_566_p2 ^ b0_11_fu_872_p3);

assign b0_80_fu_5768_p2 = (b0_84_fu_5752_p4 ^ b0_76_fu_5690_p2);

assign b0_81_fu_10457_p2 = (b0_85_reg_14510_pp0_iter1_reg ^ b0_77_fu_10170_p2);

assign b0_82_fu_10538_p2 = (b0_83_reg_14524_pp0_iter1_reg ^ b0_81_fu_10457_p2);

assign b0_84_fu_5752_p4 = {{b_274_fu_5662_p2[5:4]}};

assign b0_86_fu_10783_p2 = (b0_87_reg_14549_pp0_iter1_reg ^ b0_85_reg_14510_pp0_iter1_reg);

assign b0_88_fu_288_p4 = {{a[25:24]}};

assign b0_89_fu_11094_p2 = (a0_336_reg_14105_pp0_iter1_reg ^ a0_335_reg_13615_pp0_iter1_reg);

assign b0_8_fu_1048_p2 = (b0_9_fu_1020_p3 ^ b0_7_fu_942_p2);

assign b0_90_fu_5900_p2 = (b0_88_fu_288_p4 ^ a0_287_fu_224_p4);

assign b0_91_fu_11281_p2 = (a0_338_reg_14121_pp0_iter1_reg ^ a0_335_reg_13615_pp0_iter1_reg);

assign b0_92_fu_11361_p2 = (b0_93_reg_14580_pp0_iter1_reg ^ b0_91_fu_11281_p2);

assign b0_94_fu_11601_p2 = (a0_338_reg_14121_pp0_iter1_reg ^ a0_288_reg_13599_pp0_iter1_reg);

assign b0_9_fu_1020_p3 = b_15_fu_890_p2[32'd2];

assign b0_fu_484_p2 = (a1_258_fu_194_p4 ^ a0_289_fu_408_p1);

assign b1_100_fu_678_p3 = b_7_fu_652_p2[32'd1];

assign b1_101_fu_744_p3 = b0_1_fu_516_p2[32'd3];

assign b1_102_fu_918_p4 = {{b_15_fu_890_p2[3:2]}};

assign b1_103_fu_948_p3 = b0_6_fu_912_p2[32'd1];

assign b1_104_fu_1054_p3 = b_20_fu_1028_p2[32'd1];

assign b1_105_fu_1120_p3 = b_15_fu_890_p2[32'd3];

assign b1_106_fu_1234_p4 = {{b0_fu_484_p2[7:6]}};

assign b1_107_fu_1252_p3 = xor_ln40_1_fu_490_p2[32'd5];

assign b1_108_fu_1358_p3 = b_33_fu_1332_p2[32'd1];

assign b1_109_fu_1424_p3 = b0_fu_484_p2[32'd7];

assign b1_110_fu_1746_p4 = {{b_41_fu_1712_p2[7:4]}};

assign b1_111_fu_1778_p4 = {{b0_14_fu_1740_p2[3:2]}};

assign b1_112_fu_1808_p3 = b0_15_fu_1772_p2[32'd1];

assign b1_113_fu_1914_p3 = b_47_fu_1888_p2[32'd1];

assign b1_114_fu_1980_p3 = b0_14_fu_1740_p2[32'd3];

assign b1_115_fu_2154_p4 = {{b_55_fu_2126_p2[3:2]}};

assign b1_116_fu_2184_p3 = b0_19_fu_2148_p2[32'd1];

assign b1_117_fu_2290_p3 = b_60_fu_2264_p2[32'd1];

assign b1_118_fu_2356_p3 = b_55_fu_2126_p2[32'd3];

assign b1_119_fu_2470_p4 = {{b_41_fu_1712_p2[7:6]}};

assign b1_120_fu_2488_p3 = xor_ln33_fu_1718_p2[32'd5];

assign b1_121_fu_2594_p3 = b_73_fu_2568_p2[32'd1];

assign b1_122_fu_2660_p3 = b_41_fu_1712_p2[32'd7];

assign b1_123_fu_2870_p4 = {{a0z1_fu_440_p2[15:12]}};

assign b1_124_fu_2890_p4 = {{xor_ln70_3_fu_458_p2[11:10]}};

assign b1_125_fu_2908_p3 = xor_ln70_2_fu_452_p2[32'd9];

assign b1_126_fu_3014_p3 = b_87_fu_2988_p2[32'd1];

assign b1_127_fu_3080_p3 = xor_ln70_3_fu_458_p2[32'd11];

assign b1_128_fu_3254_p4 = {{b_95_fu_3226_p2[3:2]}};

assign b1_129_fu_3284_p3 = b0_32_fu_3248_p2[32'd1];

assign b1_130_fu_3390_p3 = b_100_fu_3364_p2[32'd1];

assign b1_131_fu_3456_p3 = b_95_fu_3226_p2[32'd3];

assign b1_132_fu_3570_p4 = {{a0z1_fu_440_p2[15:14]}};

assign b1_133_fu_3588_p3 = xor_ln70_1_fu_446_p2[32'd13];

assign b1_134_fu_3694_p3 = b_113_fu_3668_p2[32'd1];

assign b1_135_fu_3760_p3 = a0z1_fu_440_p2[32'd15];

assign b1_136_fu_5006_p4 = {{a0z1_1_fu_4978_p2[7:4]}};

assign b1_137_fu_5032_p4 = {{b0_40_fu_5000_p2[3:2]}};

assign b1_141_fu_5194_p4 = {{b_135_fu_5166_p2[3:2]}};

assign b1_145_fu_5290_p4 = {{a0z1_1_fu_4978_p2[7:6]}};

assign b1_149_fu_6894_p4 = {{a0z1_2_fu_6872_p2[3:2]}};

assign b1_150_fu_6918_p3 = b0_53_fu_6888_p2[32'd1];

assign b1_151_fu_7024_p3 = b_166_fu_6998_p2[32'd1];

assign b1_152_fu_7090_p3 = a0z1_2_fu_6872_p2[32'd3];

assign b1_153_fu_7370_p3 = a0z1_3_fu_7350_p2[32'd1];

assign b1_155_fu_5436_p4 = {{xor_ln71_3_fu_4686_p2[11:10]}};

assign b1_157_fu_5472_p4 = {{b_208_fu_5460_p2[3:2]}};

assign b1_162_fu_5534_p4 = {{a[23:20]}};

assign b1_163_fu_5544_p4 = {{a[19:18]}};

assign b1_165_fu_5590_p4 = {{b_248_fu_5578_p2[3:2]}};

assign b1_169_fu_5638_p4 = {{a[23:22]}};

assign b1_171_fu_5680_p4 = {{b_274_fu_5662_p2[7:4]}};

assign b1_172_fu_5696_p4 = {{b0_75_fu_5674_p2[3:2]}};

assign b1_176_fu_5774_p4 = {{b_288_fu_5762_p2[3:2]}};

assign b1_180_fu_5822_p4 = {{b_274_fu_5662_p2[7:6]}};

assign b1_184_fu_5870_p4 = {{a[27:26]}};

assign b1_186_fu_5906_p4 = {{b_328_fu_5894_p2[3:2]}};

assign b1_97_fu_522_p4 = {{b0_fu_484_p2[7:4]}};

assign b1_98_fu_548_p4 = {{b0_1_fu_516_p2[3:2]}};

assign b1_99_fu_572_p3 = b0_2_fu_542_p2[32'd1];

assign b1_fu_496_p4 = {{a0z1_fu_440_p2[15:8]}};

assign b_100_fu_3364_p2 = (b1_128_fu_3254_p4 ^ b0_32_fu_3248_p2);

assign b_102_fu_3410_p2 = (b1_130_fu_3390_p3 ^ b0_34_fu_3384_p2);

assign b_106_fu_3476_p2 = (b1_131_fu_3456_p3 ^ b0_35_fu_3356_p3);

assign b_111_fu_3608_p2 = (b1_133_fu_3588_p3 ^ b0_37_fu_3208_p3);

assign b_113_fu_3668_p2 = (b1_132_fu_3570_p4 ^ b0_36_fu_3216_p4);

assign b_115_fu_3714_p2 = (b1_134_fu_3694_p3 ^ b0_38_fu_3688_p2);

assign b_119_fu_3780_p2 = (b1_135_fu_3760_p3 ^ b0_39_fu_3660_p3);

assign b_125_fu_5976_p2 = (b1_138_reg_14190 ^ b0_42_reg_14181);

assign b_127_fu_5086_p2 = (b1_137_fu_5032_p4 ^ b0_41_fu_5026_p2);

assign b_129_fu_6029_p2 = (b1_139_reg_14218 ^ b0_43_fu_6014_p2);

assign b_133_fu_6072_p2 = (b1_140_reg_14231 ^ b0_44_reg_14204);

assign b_135_fu_5166_p2 = (b1_136_fu_5006_p4 ^ b0_40_fu_5000_p2);

assign b_138_fu_6171_p2 = (b1_142_reg_14261 ^ b0_46_fu_6156_p2);

assign b_13_fu_764_p2 = (b1_101_fu_744_p3 ^ b0_5_fu_644_p3);

assign b_140_fu_5242_p2 = (b1_141_fu_5194_p4 ^ b0_45_fu_5188_p2);

assign b_142_fu_6227_p2 = (b1_143_reg_14289 ^ b0_47_fu_6211_p2);

assign b_146_fu_6270_p2 = (b1_144_reg_14302 ^ b0_48_reg_14275);

assign b_151_fu_6358_p2 = (b1_146_reg_14315 ^ b0_50_reg_14246);

assign b_153_fu_5338_p2 = (b1_145_fu_5290_p4 ^ b0_49_fu_5156_p4);

assign b_155_fu_6411_p2 = (b1_147_reg_14343 ^ b0_51_fu_6396_p2);

assign b_159_fu_6454_p2 = (b1_148_reg_14356 ^ b0_52_reg_14329);

assign b_15_fu_890_p2 = (b1_97_fu_522_p4 ^ b0_1_fu_516_p2);

assign b_164_fu_6938_p2 = (b1_150_fu_6918_p3 ^ b0_54_fu_6912_p2);

assign b_166_fu_6998_p2 = (b1_149_fu_6894_p4 ^ b0_53_fu_6888_p2);

assign b_168_fu_7044_p2 = (b1_151_fu_7024_p3 ^ b0_55_fu_7018_p2);

assign b_172_fu_7110_p2 = (b1_152_fu_7090_p3 ^ b0_56_fu_6990_p3);

assign b_176_fu_7390_p2 = (b1_153_fu_7370_p3 ^ b0_57_fu_7356_p2);

assign b_181_fu_7336_p2 = (a1_343_fu_7328_p3 ^ a0_372_fu_7320_p3);

assign b_185_fu_7222_p2 = (a1_342_fu_7214_p3 ^ a0_369_fu_7206_p3);

assign b_187_fu_7558_p2 = (a1_336_fu_6759_p4 ^ a0_363_fu_6749_p4);

assign b_189_fu_7656_p2 = (b1_154_reg_14798 ^ b0_58_fu_7640_p2);

assign b_18_fu_968_p2 = (b1_103_fu_948_p3 ^ b0_7_fu_942_p2);

assign b_198_fu_6624_p2 = (a1_333_reg_14371 ^ a0_357_reg_14363);

assign b_200_fu_5446_p2 = (b1_155_fu_5436_p4 ^ b0_59_fu_4800_p4);

assign b_202_fu_7998_p2 = (b1_156_reg_14411_pp0_iter1_reg ^ b0_60_fu_7982_p2);

assign b_208_fu_5460_p2 = (a1_316_fu_4726_p4 ^ a0_341_fu_4716_p4);

assign b_20_fu_1028_p2 = (b1_102_fu_918_p4 ^ b0_6_fu_912_p2);

assign b_211_fu_8185_p2 = (b1_158_reg_14417_pp0_iter1_reg ^ b0_62_fu_8169_p2);

assign b_213_fu_5498_p2 = (b1_157_fu_5472_p4 ^ b0_61_fu_5466_p2);

assign b_215_fu_8266_p2 = (b1_159_reg_14430_pp0_iter1_reg ^ b0_63_fu_8249_p2);

assign b_219_fu_8321_p2 = (b1_160_reg_14436_pp0_iter1_reg ^ b0_64_reg_14423_pp0_iter1_reg);

assign b_224_fu_6659_p2 = (a1_335_reg_14397 ^ a0_360_reg_14159);

assign b_226_fu_5520_p2 = (a1_317_fu_4746_p4 ^ a0_342_fu_4736_p4);

assign b_228_fu_8491_p2 = (b1_161_reg_14442_pp0_iter1_reg ^ b0_65_fu_8475_p2);

assign b_22_fu_1074_p2 = (b1_104_fu_1054_p3 ^ b0_8_fu_1048_p2);

assign b_238_fu_4172_p2 = (a1_307_fu_4164_p3 ^ a0_329_fu_4156_p3);

assign b_240_fu_5554_p2 = (b1_163_fu_5544_p4 ^ b0_67_fu_328_p4);

assign b_242_fu_9384_p2 = (b1_164_reg_14448_pp0_iter1_reg ^ b0_68_fu_9368_p2);

assign b_248_fu_5578_p2 = (b1_162_fu_5534_p4 ^ b0_66_fu_318_p4);

assign b_251_fu_9569_p2 = (b1_166_reg_14454_pp0_iter1_reg ^ b0_70_fu_9553_p2);

assign b_253_fu_5616_p2 = (b1_165_fu_5590_p4 ^ b0_69_fu_5584_p2);

assign b_255_fu_9650_p2 = (b1_167_reg_14467_pp0_iter1_reg ^ b0_71_fu_9633_p2);

assign b_259_fu_9705_p2 = (b1_168_reg_14473_pp0_iter1_reg ^ b0_72_reg_14460_pp0_iter1_reg);

assign b_264_fu_4256_p2 = (a1_309_fu_4248_p3 ^ a0_332_fu_4240_p3);

assign b_266_fu_5648_p2 = (b1_169_fu_5638_p4 ^ b0_73_fu_5568_p4);

assign b_268_fu_9889_p2 = (b1_170_reg_14479_pp0_iter1_reg ^ b0_74_fu_9873_p2);

assign b_26_fu_1140_p2 = (b1_105_fu_1120_p3 ^ b0_9_fu_1020_p3);

assign b_274_fu_5662_p2 = (a1_258_fu_194_p4 ^ a0_285_fu_184_p4);

assign b_278_fu_10186_p2 = (b1_173_reg_14485_pp0_iter1_reg ^ b0_77_fu_10170_p2);

assign b_280_fu_5722_p2 = (b1_172_fu_5696_p4 ^ b0_76_fu_5690_p2);

assign b_282_fu_10267_p2 = (b1_174_reg_14498_pp0_iter1_reg ^ b0_78_fu_10250_p2);

assign b_286_fu_10322_p2 = (b1_175_reg_14504_pp0_iter1_reg ^ b0_79_reg_14491_pp0_iter1_reg);

assign b_288_fu_5762_p2 = (b1_171_fu_5680_p4 ^ b0_75_fu_5674_p2);

assign b_291_fu_10474_p2 = (b1_177_reg_14518_pp0_iter1_reg ^ b0_81_fu_10457_p2);

assign b_293_fu_5800_p2 = (b1_176_fu_5774_p4 ^ b0_80_fu_5768_p2);

assign b_295_fu_10555_p2 = (b1_178_reg_14531_pp0_iter1_reg ^ b0_82_fu_10538_p2);

assign b_299_fu_10610_p2 = (b1_179_reg_14537_pp0_iter1_reg ^ b0_83_reg_14524_pp0_iter1_reg);

assign b_304_fu_10720_p2 = (b1_181_reg_14543_pp0_iter1_reg ^ b0_85_reg_14510_pp0_iter1_reg);

assign b_306_fu_5848_p2 = (b1_180_fu_5822_p4 ^ b0_84_fu_5752_p4);

assign b_308_fu_10799_p2 = (b1_182_reg_14556_pp0_iter1_reg ^ b0_86_fu_10783_p2);

assign b_312_fu_10854_p2 = (b1_183_reg_14562_pp0_iter1_reg ^ b0_87_reg_14549_pp0_iter1_reg);

assign b_318_fu_4362_p2 = (a1_311_fu_4354_p3 ^ a0_335_fu_362_p3);

assign b_31_fu_1272_p2 = (b1_107_fu_1252_p3 ^ b0_11_fu_872_p3);

assign b_320_fu_5880_p2 = (b1_184_fu_5870_p4 ^ b0_88_fu_288_p4);

assign b_322_fu_11110_p2 = (b1_185_reg_14568_pp0_iter1_reg ^ b0_89_fu_11094_p2);

assign b_328_fu_5894_p2 = (a1_259_fu_214_p4 ^ a0_286_fu_204_p4);

assign b_331_fu_11297_p2 = (b1_187_reg_14574_pp0_iter1_reg ^ b0_91_fu_11281_p2);

assign b_333_fu_5932_p2 = (b1_186_fu_5906_p4 ^ b0_90_fu_5900_p2);

assign b_335_fu_11378_p2 = (b1_188_reg_14587_pp0_iter1_reg ^ b0_92_fu_11361_p2);

assign b_339_fu_11433_p2 = (b1_189_reg_14593_pp0_iter1_reg ^ b0_93_reg_14580_pp0_iter1_reg);

assign b_33_fu_1332_p2 = (b1_106_fu_1234_p4 ^ b0_10_fu_880_p4);

assign b_344_fu_4446_p2 = (a1_313_fu_4438_p3 ^ a0_338_fu_4430_p3);

assign b_346_fu_5954_p2 = (a1_260_fu_234_p4 ^ a0_287_fu_224_p4);

assign b_348_fu_11617_p2 = (b1_190_reg_14599_pp0_iter1_reg ^ b0_94_fu_11601_p2);

assign b_35_fu_1378_p2 = (b1_108_fu_1358_p3 ^ b0_12_fu_1352_p2);

assign b_39_fu_1444_p2 = (b1_109_fu_1424_p3 ^ b0_13_fu_1324_p3);

assign b_41_fu_1712_p2 = (b1_fu_496_p4 ^ b0_fu_484_p2);

assign b_45_fu_1828_p2 = (b1_112_fu_1808_p3 ^ b0_16_fu_1802_p2);

assign b_47_fu_1888_p2 = (b1_111_fu_1778_p4 ^ b0_15_fu_1772_p2);

assign b_49_fu_1934_p2 = (b1_113_fu_1914_p3 ^ b0_17_fu_1908_p2);

assign b_53_fu_2000_p2 = (b1_114_fu_1980_p3 ^ b0_18_fu_1880_p3);

assign b_55_fu_2126_p2 = (b1_110_fu_1746_p4 ^ b0_14_fu_1740_p2);

assign b_58_fu_2204_p2 = (b1_116_fu_2184_p3 ^ b0_20_fu_2178_p2);

assign b_5_fu_592_p2 = (b1_99_fu_572_p3 ^ b0_3_fu_566_p2);

assign b_60_fu_2264_p2 = (b1_115_fu_2154_p4 ^ b0_19_fu_2148_p2);

assign b_62_fu_2310_p2 = (b1_117_fu_2290_p3 ^ b0_21_fu_2284_p2);

assign b_66_fu_2376_p2 = (b1_118_fu_2356_p3 ^ b0_22_fu_2256_p3);

assign b_71_fu_2508_p2 = (b1_120_fu_2488_p3 ^ b0_24_fu_2108_p3);

assign b_73_fu_2568_p2 = (b1_119_fu_2470_p4 ^ b0_23_fu_2116_p4);

assign b_75_fu_2614_p2 = (b1_121_fu_2594_p3 ^ b0_25_fu_2588_p2);

assign b_79_fu_2680_p2 = (b1_122_fu_2660_p3 ^ b0_26_fu_2560_p3);

assign b_7_fu_652_p2 = (b1_98_fu_548_p4 ^ b0_2_fu_542_p2);

assign b_85_fu_2928_p2 = (b1_125_fu_2908_p3 ^ b0_29_fu_1674_p3);

assign b_87_fu_2988_p2 = (b1_124_fu_2890_p4 ^ b0_28_fu_1682_p4);

assign b_89_fu_3034_p2 = (b1_126_fu_3014_p3 ^ b0_30_fu_3008_p2);

assign b_93_fu_3100_p2 = (b1_127_fu_3080_p3 ^ b0_31_fu_2980_p3);

assign b_95_fu_3226_p2 = (b1_123_fu_2870_p4 ^ b0_27_fu_1692_p4);

assign b_98_fu_3304_p2 = (b1_129_fu_3284_p3 ^ b0_33_fu_3278_p2);

assign b_9_fu_698_p2 = (b1_100_fu_678_p3 ^ b0_4_fu_672_p2);

assign delta_1_fu_6731_p2 = (tmp_37_fu_6707_p4 ^ tmp_35_fu_6616_p3);

assign delta_2_fu_7284_p2 = (tmp_42_fu_7260_p3 ^ tmp_41_fu_7198_p3);

assign delta_3_fu_7436_p2 = (tmp_45_fu_7428_p3 ^ tmp_44_fu_7420_p3);

assign delta_4_fu_7468_p2 = (and_ln36_fu_7462_p2 ^ a1_345_fu_7448_p3);

assign delta_fu_4668_p2 = (tmp_26_fu_4602_p5 ^ tmp_21_fu_4148_p3);

assign tmp_100_fu_4046_p3 = {{xor_ln45_85_fu_2846_p2}, {xor_ln45_67_fu_2834_p2}};

assign tmp_101_fu_4060_p3 = {{xor_ln28_28_fu_4024_p2}, {a1_305_fu_3928_p2}};

assign tmp_102_fu_4068_p3 = {{xor_ln45_130_fu_3940_p2}, {a0_73_fu_3934_p2}};

assign tmp_103_fu_4574_p3 = {{tmp_213_fu_4306_p4}, {xor_ln59_6_fu_4338_p2}};

assign tmp_104_fu_4582_p3 = {{a1_314_fu_4474_p4}, {a0_96_fu_4506_p2}};

assign tmp_105_fu_4614_p3 = {{xor_ln45_152_fu_4142_p2}, {xor_ln45_105_fu_4124_p2}};

assign tmp_106_fu_4622_p4 = {{{a1_315_fu_4500_p2}, {a1_314_fu_4474_p4}}, {xor_ln59_13_fu_4590_p2}};

assign tmp_107_fu_4632_p3 = {{xor_ln45_147_fu_4136_p2}, {xor_ln45_105_fu_4124_p2}};

assign tmp_108_fu_4640_p3 = {{a1_314_fu_4474_p4}, {xor_ln59_13_fu_4590_p2}};

assign tmp_109_fu_4648_p3 = {{xor_ln45_146_fu_4130_p2}, {xor_ln45_105_fu_4124_p2}};

assign tmp_10_fu_2724_p3 = {{xor_ln28_11_fu_2718_p2}, {a1_46_fu_2698_p2}};

assign tmp_110_fu_4656_p5 = {{{{xor_ln59_14_fu_4596_p2}, {a1_315_fu_4500_p2}}, {a1_314_fu_4474_p4}}, {xor_ln59_13_fu_4590_p2}};

assign tmp_111_fu_4970_p3 = {{xor_ln28_42_fu_4824_p2}, {a1_316_fu_4726_p4}};

assign tmp_112_fu_6716_p3 = {{xor_ln45_183_fu_6610_p2}, {xor_ln45_139_fu_6604_p2}};

assign tmp_113_fu_6724_p3 = {{tmp_258_reg_14404}, {xor_ln59_19_fu_6701_p2}};

assign tmp_114_fu_7268_p3 = {{xor_ln45_201_fu_7192_p2}, {xor_ln45_149_fu_7186_p2}};

assign tmp_115_fu_7276_p3 = {{a1_337_fu_6777_p3}, {xor_ln59_21_fu_7244_p2}};

assign tmp_11_fu_2782_p3 = {{xor_ln28_12_fu_2776_p2}, {a1_49_fu_2768_p3}};

assign tmp_12_fu_2796_p3 = {{xor_ln28_13_fu_2790_p2}, {a1_290_fu_2744_p2}};

assign tmp_13_fu_3144_p3 = {{xor_ln28_14_fu_3138_p2}, {a1_56_fu_3118_p2}};

assign tmp_14_fu_3520_p3 = {{xor_ln28_15_fu_3514_p2}, {a1_61_fu_3494_p2}};

assign tmp_15_fu_3824_p3 = {{xor_ln28_16_fu_3818_p2}, {a1_66_fu_3798_p2}};

assign tmp_16_fu_3882_p3 = {{xor_ln28_17_fu_3876_p2}, {a1_68_fu_3868_p3}};

assign tmp_17_fu_3896_p3 = {{xor_ln28_18_fu_3890_p2}, {a1_304_fu_3844_p2}};

assign tmp_18_fu_3996_p3 = {{xor_ln28_19_fu_3990_p2}, {a1_71_fu_3982_p3}};

assign tmp_19_fu_4010_p3 = {{xor_ln28_20_fu_4004_p2}, {a1_306_fu_3964_p4}};

assign tmp_1_fu_280_p3 = {{xor_ln28_1_fu_274_p2}, {a1_260_fu_234_p4}};

integer ap_tvar_int_1;

always @ (a) begin
    for (ap_tvar_int_1 = 2 - 1; ap_tvar_int_1 >= 0; ap_tvar_int_1 = ap_tvar_int_1 - 1) begin
        if (ap_tvar_int_1 > 19 - 18) begin
            tmp_208_fu_4222_p4[ap_tvar_int_1] = 1'b0;
        end else begin
            tmp_208_fu_4222_p4[ap_tvar_int_1] = a[19 - ap_tvar_int_1];
        end
    end
end

assign tmp_20_fu_4030_p3 = {{xor_ln28_21_fu_4018_p2}, {a1_305_fu_3928_p2}};

integer ap_tvar_int_2;

always @ (a) begin
    for (ap_tvar_int_2 = 2 - 1; ap_tvar_int_2 >= 0; ap_tvar_int_2 = ap_tvar_int_2 - 1) begin
        if (ap_tvar_int_2 > 23 - 22) begin
            tmp_213_fu_4306_p4[ap_tvar_int_2] = 1'b0;
        end else begin
            tmp_213_fu_4306_p4[ap_tvar_int_2] = a[23 - ap_tvar_int_2];
        end
    end
end

integer ap_tvar_int_3;

always @ (a) begin
    for (ap_tvar_int_3 = 2 - 1; ap_tvar_int_3 >= 0; ap_tvar_int_3 = ap_tvar_int_3 - 1) begin
        if (ap_tvar_int_3 > 27 - 26) begin
            tmp_217_fu_4412_p4[ap_tvar_int_3] = 1'b0;
        end else begin
            tmp_217_fu_4412_p4[ap_tvar_int_3] = a[27 - ap_tvar_int_3];
        end
    end
end

assign tmp_21_fu_4148_p3 = {{xor_ln45_104_fu_4118_p2}, {xor_ln45_105_fu_4124_p2}};

assign tmp_22_fu_4324_p3 = {{a0_334_fu_4286_p2}, {a0_333_fu_4270_p3}};

assign tmp_23_fu_4492_p3 = {{a0_339_fu_260_p2}, {a0_288_fu_244_p3}};

assign tmp_24_fu_4540_p3 = {{xor_ln28_30_fu_4534_p2}, {a1_88_fu_4526_p3}};

integer ap_tvar_int_4;

always @ (xor_ln71_3_fu_4686_p2) begin
    for (ap_tvar_int_4 = 2 - 1; ap_tvar_int_4 >= 0; ap_tvar_int_4 = ap_tvar_int_4 - 1) begin
        if (ap_tvar_int_4 > 11 - 10) begin
            tmp_256_fu_5408_p4[ap_tvar_int_4] = 1'b0;
        end else begin
            tmp_256_fu_5408_p4[ap_tvar_int_4] = xor_ln71_3_fu_4686_p2[11 - ap_tvar_int_4];
        end
    end
end

integer ap_tvar_int_5;

always @ (delta_fu_4668_p2) begin
    for (ap_tvar_int_5 = 2 - 1; ap_tvar_int_5 >= 0; ap_tvar_int_5 = ap_tvar_int_5 - 1) begin
        if (ap_tvar_int_5 > 15 - 14) begin
            tmp_258_fu_5426_p4[ap_tvar_int_5] = 1'b0;
        end else begin
            tmp_258_fu_5426_p4[ap_tvar_int_5] = delta_fu_4668_p2[15 - ap_tvar_int_5];
        end
    end
end

assign tmp_25_fu_4554_p3 = {{xor_ln28_31_fu_4548_p2}, {a1_315_fu_4500_p2}};

assign tmp_26_fu_4602_p5 = {{{{xor_ln28_32_fu_4568_p2}, {a1_315_fu_4500_p2}}, {a1_314_fu_4474_p4}}, {xor_ln59_13_fu_4590_p2}};

integer ap_tvar_int_6;

always @ (delta_1_fu_6731_p2) begin
    for (ap_tvar_int_6 = 2 - 1; ap_tvar_int_6 >= 0; ap_tvar_int_6 = ap_tvar_int_6 - 1) begin
        if (ap_tvar_int_6 > 7 - 6) begin
            tmp_271_fu_7250_p4[ap_tvar_int_6] = 1'b0;
        end else begin
            tmp_271_fu_7250_p4[ap_tvar_int_6] = delta_1_fu_6731_p2[7 - ap_tvar_int_6];
        end
    end
end

assign tmp_27_fu_4778_p3 = {{a0_361_fu_4772_p2}, {a1_318_fu_4764_p3}};

assign tmp_28_fu_4792_p3 = {{xor_ln28_34_fu_4786_p2}, {a1_317_fu_4746_p4}};

assign tmp_29_fu_4830_p3 = {{xor_ln28_35_fu_4810_p2}, {a1_316_fu_4726_p4}};

assign tmp_2_fu_310_p3 = {{xor_ln28_2_fu_298_p2}, {a1_259_fu_214_p4}};

assign tmp_30_fu_6112_p3 = {{xor_ln28_36_fu_6106_p2}, {a1_98_fu_6086_p2}};

assign tmp_31_fu_6310_p3 = {{xor_ln28_37_fu_6304_p2}, {a1_103_fu_6284_p2}};

assign tmp_32_fu_6494_p3 = {{xor_ln28_38_fu_6488_p2}, {a1_109_fu_6468_p2}};

assign tmp_33_fu_6552_p3 = {{xor_ln28_39_fu_6546_p2}, {a1_111_fu_6538_p3}};

assign tmp_34_fu_6566_p3 = {{xor_ln28_40_fu_6560_p2}, {a1_332_fu_6514_p2}};

assign tmp_35_fu_6616_p3 = {{xor_ln45_138_fu_6598_p2}, {xor_ln45_139_fu_6604_p2}};

assign tmp_36_fu_6689_p3 = {{a0_361_reg_14151}, {a0_343_reg_14138}};

assign tmp_37_fu_6707_p4 = {{{xor_ln28_43_fu_6695_p2}, {tmp_258_reg_14404}}, {xor_ln59_19_fu_6701_p2}};

assign tmp_38_fu_6791_p3 = {{a0_370_fu_6785_p2}, {a1_337_fu_6777_p3}};

assign tmp_39_fu_6805_p3 = {{xor_ln28_45_fu_6799_p2}, {a1_336_fu_6759_p4}};

assign tmp_3_fu_388_p3 = {{xor_ln28_3_fu_356_p2}, {a1_258_fu_194_p4}};

assign tmp_40_fu_7154_p3 = {{xor_ln28_46_fu_7148_p2}, {a1_126_fu_7128_p2}};

assign tmp_41_fu_7198_p3 = {{xor_ln45_148_fu_7180_p2}, {xor_ln45_149_fu_7186_p2}};

assign tmp_42_fu_7260_p3 = {{tmp_271_fu_7250_p4}, {xor_ln59_21_fu_7244_p2}};

assign tmp_43_fu_7342_p3 = {{b_181_fu_7336_p2}, {a1_343_fu_7328_p3}};

assign tmp_44_fu_7420_p3 = {{xor_ln45_150_fu_7408_p2}, {xor_ln45_151_fu_7414_p2}};

assign tmp_45_fu_7428_p3 = {{a1_343_fu_7328_p3}, {b_181_fu_7336_p2}};

assign tmp_46_fu_7730_p3 = {{xor_ln28_48_fu_7724_p2}, {a1_141_fu_7704_p2}};

assign tmp_47_fu_7867_p3 = {{xor_ln28_49_fu_7861_p2}, {a1_142_fu_7841_p2}};

assign tmp_48_fu_8089_p3 = {{xor_ln28_50_fu_8083_p2}, {a1_149_fu_8063_p2}};

assign tmp_49_fu_8362_p3 = {{xor_ln28_51_fu_8356_p2}, {a1_155_fu_8336_p2}};

assign tmp_4_fu_1488_p3 = {{xor_ln28_6_fu_1482_p2}, {a1_24_fu_1462_p2}};

assign tmp_50_fu_8582_p3 = {{xor_ln28_52_fu_8576_p2}, {a1_161_fu_8556_p2}};

assign tmp_51_fu_8640_p3 = {{xor_ln28_53_fu_8634_p2}, {a1_163_fu_8626_p3}};

assign tmp_52_fu_8654_p3 = {{xor_ln28_54_fu_8648_p2}, {a1_364_fu_8602_p2}};

assign tmp_53_fu_8809_p3 = {{xor_ln28_55_fu_8803_p2}, {a1_164_fu_8783_p2}};

assign tmp_54_fu_8960_p3 = {{xor_ln28_56_fu_8954_p2}, {a1_165_fu_8934_p2}};

assign tmp_55_fu_9111_p3 = {{xor_ln28_57_fu_9105_p2}, {a1_167_fu_9085_p2}};

assign tmp_56_fu_9169_p3 = {{xor_ln28_58_fu_9163_p2}, {a1_169_fu_9155_p3}};

assign tmp_57_fu_9183_p3 = {{xor_ln28_59_fu_9177_p2}, {a1_365_fu_9131_p2}};

assign tmp_58_fu_9475_p3 = {{xor_ln28_60_fu_9469_p2}, {a1_178_fu_9449_p2}};

assign tmp_59_fu_9746_p3 = {{xor_ln28_61_fu_9740_p2}, {a1_183_fu_9720_p2}};

assign tmp_5_fu_1546_p3 = {{xor_ln28_7_fu_1540_p2}, {a1_27_fu_1532_p3}};

assign tmp_60_fu_9980_p3 = {{xor_ln28_62_fu_9974_p2}, {a1_190_fu_9954_p2}};

assign tmp_61_fu_10038_p3 = {{xor_ln28_63_fu_10032_p2}, {a1_192_fu_10024_p3}};

assign tmp_62_fu_10052_p3 = {{xor_ln28_64_fu_10046_p2}, {a1_380_fu_10000_p2}};

assign tmp_63_fu_10363_p3 = {{xor_ln28_65_fu_10357_p2}, {a1_198_fu_10337_p2}};

assign tmp_64_fu_10651_p3 = {{xor_ln28_66_fu_10645_p2}, {a1_212_fu_10625_p2}};

assign tmp_65_fu_10895_p3 = {{xor_ln28_67_fu_10889_p2}, {a1_217_fu_10869_p2}};

assign tmp_66_fu_10953_p3 = {{xor_ln28_68_fu_10947_p2}, {a1_219_fu_10939_p3}};

assign tmp_67_fu_10967_p3 = {{xor_ln28_69_fu_10961_p2}, {a1_394_fu_10915_p2}};

assign tmp_68_fu_11201_p3 = {{xor_ln28_70_fu_11195_p2}, {a1_225_fu_11175_p2}};

assign tmp_69_fu_11474_p3 = {{xor_ln28_71_fu_11468_p2}, {a1_230_fu_11448_p2}};

assign tmp_6_fu_1560_p3 = {{xor_ln28_8_fu_1554_p2}, {a1_276_fu_1508_p2}};

assign tmp_70_fu_11708_p3 = {{xor_ln28_fu_11702_p2}, {a1_fu_11682_p2}};

assign tmp_71_fu_11766_p3 = {{xor_ln28_72_fu_11760_p2}, {a1_236_fu_11752_p3}};

assign tmp_72_fu_11780_p3 = {{xor_ln28_73_fu_11774_p2}, {a1_408_fu_11728_p2}};

assign tmp_73_fu_11856_p3 = {{xor_ln28_74_fu_11850_p2}, {a1_239_fu_11842_p3}};

assign tmp_74_fu_11870_p3 = {{xor_ln28_75_fu_11864_p2}, {a1_410_fu_11824_p4}};

assign tmp_75_fu_11884_p3 = {{xor_ln28_76_fu_11878_p2}, {a1_409_fu_11800_p2}};

assign tmp_76_fu_12027_p3 = {{xor_ln28_77_fu_12021_p2}, {a1_240_fu_12001_p2}};

assign tmp_77_fu_12178_p3 = {{xor_ln28_78_fu_12172_p2}, {a1_241_fu_12152_p2}};

assign tmp_78_fu_12329_p3 = {{xor_ln28_79_fu_12323_p2}, {a1_242_fu_12303_p2}};

assign tmp_79_fu_12387_p3 = {{xor_ln28_80_fu_12381_p2}, {a1_244_fu_12373_p3}};

assign tmp_7_fu_808_p3 = {{xor_ln28_4_fu_802_p2}, {a1_13_fu_782_p2}};

assign tmp_80_fu_12401_p3 = {{xor_ln28_81_fu_12395_p2}, {a1_411_fu_12349_p2}};

assign tmp_81_fu_12552_p3 = {{xor_ln28_82_fu_12546_p2}, {a1_245_fu_12526_p2}};

assign tmp_82_fu_12703_p3 = {{xor_ln28_83_fu_12697_p2}, {a1_246_fu_12677_p2}};

assign tmp_83_fu_12854_p3 = {{xor_ln28_84_fu_12848_p2}, {a1_247_fu_12828_p2}};

assign tmp_84_fu_12912_p3 = {{xor_ln28_85_fu_12906_p2}, {a1_249_fu_12898_p3}};

assign tmp_85_fu_12926_p3 = {{xor_ln28_86_fu_12920_p2}, {a1_412_fu_12874_p2}};

assign tmp_86_fu_13077_p3 = {{xor_ln28_87_fu_13071_p2}, {a1_250_fu_13051_p2}};

assign tmp_87_fu_13228_p3 = {{xor_ln28_88_fu_13222_p2}, {a1_251_fu_13202_p2}};

assign tmp_88_fu_13379_p3 = {{xor_ln28_89_fu_13373_p2}, {a1_252_fu_13353_p2}};

assign tmp_89_fu_13437_p3 = {{xor_ln28_90_fu_13431_p2}, {a1_254_fu_13423_p3}};

assign tmp_8_fu_2044_p3 = {{xor_ln28_9_fu_2038_p2}, {a1_34_fu_2018_p2}};

assign tmp_90_fu_13451_p3 = {{xor_ln28_91_fu_13445_p2}, {a1_413_fu_13399_p2}};

assign tmp_91_fu_13527_p3 = {{xor_ln28_92_fu_13521_p2}, {a1_257_fu_13513_p3}};

assign tmp_92_fu_13541_p3 = {{xor_ln28_93_fu_13535_p2}, {a1_415_fu_13495_p4}};

assign tmp_93_fu_13555_p3 = {{xor_ln28_94_fu_13549_p2}, {a1_414_fu_13471_p2}};

assign tmp_95_fu_348_p3 = {{xor_ln28_23_fu_304_p2}, {a1_259_fu_214_p4}};

assign tmp_96_fu_416_p3 = {{xor_ln28_27_fu_382_p2}, {a1_258_fu_194_p4}};

assign tmp_97_fu_424_p3 = {{xor_ln28_26_fu_376_p2}, {a1_258_fu_194_p4}};

assign tmp_98_fu_432_p3 = {{xor_ln28_24_fu_370_p2}, {a1_258_fu_194_p4}};

assign tmp_99_fu_4038_p3 = {{xor_ln45_40_fu_1604_p2}, {xor_ln45_33_fu_1598_p2}};

assign tmp_9_fu_2420_p3 = {{xor_ln28_10_fu_2414_p2}, {a1_40_fu_2394_p2}};

assign tmp_fu_266_p3 = {{a0_339_fu_260_p2}, {a1_261_fu_252_p3}};

assign tmp_s_fu_1184_p3 = {{xor_ln28_5_fu_1178_p2}, {a1_19_fu_1158_p2}};

assign trunc_ln28_4_fu_338_p4 = {{a[21:16]}};

assign trunc_ln40_1_fu_474_p4 = {{a[29:24]}};

assign trunc_ln43_1_fu_1702_p4 = {{a0z1_fu_440_p2[13:8]}};

assign trunc_ln43_2_fu_10104_p3 = {{a0_429_fu_10100_p1}, {a0_420_fu_8692_p2}};

assign trunc_ln43_s_fu_1652_p4 = {{a[13:8]}};

assign trunc_ln68_1_fu_172_p1 = a[13:0];

assign trunc_ln68_2_fu_176_p1 = a[9:0];

assign trunc_ln68_3_fu_180_p1 = a[11:0];

assign trunc_ln70_4_fu_412_p1 = a[5:0];

assign xor_ln28_10_fu_2414_p2 = (z2_19_fu_2388_p2 ^ z1_20_fu_2382_p2);

assign xor_ln28_11_fu_2718_p2 = (z2_23_fu_2692_p2 ^ z1_25_fu_2686_p2);

assign xor_ln28_12_fu_2776_p2 = (a1_49_fu_2768_p3 ^ a0_52_fu_2764_p1);

assign xor_ln28_13_fu_2790_p2 = (tmp_11_fu_2782_p3 ^ a0_50_fu_2750_p2);

assign xor_ln28_14_fu_3138_p2 = (z2_28_fu_3112_p2 ^ z1_30_fu_3106_p2);

assign xor_ln28_15_fu_3514_p2 = (z2_32_fu_3488_p2 ^ z1_34_fu_3482_p2);

assign xor_ln28_16_fu_3818_p2 = (z2_36_fu_3792_p2 ^ z1_39_fu_3786_p2);

assign xor_ln28_17_fu_3876_p2 = (a1_68_fu_3868_p3 ^ a0_72_fu_3864_p1);

assign xor_ln28_18_fu_3890_p2 = (tmp_16_fu_3882_p3 ^ a0_70_fu_3850_p2);

assign xor_ln28_19_fu_3990_p2 = (a1_71_fu_3982_p3 ^ a0_76_fu_3974_p3);

assign xor_ln28_1_fu_274_p2 = (tmp_fu_266_p3 ^ a0_287_fu_224_p4);

assign xor_ln28_20_fu_4004_p2 = (tmp_18_fu_3996_p3 ^ a0_74_fu_3960_p1);

assign xor_ln28_21_fu_4018_p2 = (tmp_19_fu_4010_p3 ^ a0_73_fu_3934_p2);

assign xor_ln28_23_fu_304_p2 = (b0_88_fu_288_p4 ^ a1_260_fu_234_p4);

assign xor_ln28_24_fu_370_p2 = (trunc_ln28_4_fu_338_p4 ^ tmp_95_fu_348_p3);

assign xor_ln28_25_fu_4332_p2 = (tmp_22_fu_4324_p3 ^ a0_86_fu_4300_p2);

assign xor_ln28_26_fu_376_p2 = (b0_67_fu_328_p4 ^ a0_287_fu_224_p4);

assign xor_ln28_27_fu_382_p2 = (b0_66_fu_318_p4 ^ a1_259_fu_214_p4);

assign xor_ln28_28_fu_4024_p2 = (xor_ln45_131_fu_3946_p2 ^ a1_306_fu_3964_p4);

assign xor_ln28_2_fu_298_p2 = (tmp_1_fu_280_p3 ^ a0_286_fu_204_p4);

assign xor_ln28_30_fu_4534_p2 = (a1_88_fu_4526_p3 ^ a0_98_fu_4522_p1);

assign xor_ln28_31_fu_4548_p2 = (tmp_24_fu_4540_p3 ^ a1_314_fu_4474_p4);

assign xor_ln28_32_fu_4568_p2 = (tmp_25_fu_4554_p3 ^ a0_96_fu_4506_p2);

assign xor_ln28_33_fu_4562_p2 = (xor_ln59_9_fu_4406_p2 ^ a0_94_fu_4468_p2);

assign xor_ln28_34_fu_4786_p2 = (tmp_27_fu_4778_p3 ^ a0_342_fu_4736_p4);

assign xor_ln28_35_fu_4810_p2 = (tmp_28_fu_4792_p3 ^ a0_341_fu_4716_p4);

assign xor_ln28_36_fu_6106_p2 = (z2_42_fu_6082_p2 ^ z1_43_fu_6076_p2);

assign xor_ln28_37_fu_6304_p2 = (z2_46_fu_6280_p2 ^ z1_47_fu_6274_p2);

assign xor_ln28_38_fu_6488_p2 = (z2_50_fu_6464_p2 ^ z1_52_fu_6458_p2);

assign xor_ln28_39_fu_6546_p2 = (a1_111_fu_6538_p3 ^ a0_130_fu_6534_p1);

assign xor_ln28_3_fu_356_p2 = (tmp_2_fu_310_p3 ^ a0_285_fu_184_p4);

assign xor_ln28_40_fu_6560_p2 = (tmp_33_fu_6552_p3 ^ a0_129_fu_6520_p2);

assign xor_ln28_42_fu_4824_p2 = (b0_59_fu_4800_p4 ^ a1_317_fu_4746_p4);

assign xor_ln28_43_fu_6695_p2 = (tmp_36_fu_6689_p3 ^ a0_138_fu_6676_p2);

assign xor_ln28_45_fu_6799_p2 = (tmp_38_fu_6791_p3 ^ a0_363_fu_6749_p4);

assign xor_ln28_46_fu_7148_p2 = (z2_55_fu_7122_p2 ^ z1_56_fu_7116_p2);

assign xor_ln28_48_fu_7724_p2 = (z2_62_fu_7700_p2 ^ z1_63_fu_7696_p2);

assign xor_ln28_49_fu_7861_p2 = (z2_66_fu_7837_p2 ^ z1_67_fu_7833_p2);

assign xor_ln28_4_fu_802_p2 = (z2_2_fu_776_p2 ^ z1_3_fu_770_p2);

assign xor_ln28_50_fu_8083_p2 = (z2_70_fu_8058_p2 ^ z1_71_fu_8053_p2);

assign xor_ln28_51_fu_8356_p2 = (z2_74_fu_8331_p2 ^ z1_75_fu_8325_p2);

assign xor_ln28_52_fu_8576_p2 = (z2_78_fu_8551_p2 ^ z1_80_fu_8546_p2);

assign xor_ln28_53_fu_8634_p2 = (a1_163_fu_8626_p3 ^ a0_202_fu_8622_p1);

assign xor_ln28_54_fu_8648_p2 = (tmp_51_fu_8640_p3 ^ a0_201_fu_8608_p2);

assign xor_ln28_55_fu_8803_p2 = (z2_83_fu_8778_p2 ^ z1_84_fu_8773_p2);

assign xor_ln28_56_fu_8954_p2 = (z2_87_fu_8929_p2 ^ z1_88_fu_8924_p2);

assign xor_ln28_57_fu_9105_p2 = (z2_91_fu_9080_p2 ^ z1_93_fu_9075_p2);

assign xor_ln28_58_fu_9163_p2 = (a1_169_fu_9155_p3 ^ a0_207_fu_9151_p1);

assign xor_ln28_59_fu_9177_p2 = (tmp_56_fu_9169_p3 ^ a0_206_fu_9137_p2);

assign xor_ln28_5_fu_1178_p2 = (z2_6_fu_1152_p2 ^ z1_7_fu_1146_p2);

assign xor_ln28_60_fu_9469_p2 = (z2_96_fu_9444_p2 ^ z1_97_fu_9439_p2);

assign xor_ln28_61_fu_9740_p2 = (z2_100_fu_9715_p2 ^ z1_101_fu_9709_p2);

assign xor_ln28_62_fu_9974_p2 = (z2_104_fu_9949_p2 ^ z1_106_fu_9944_p2);

assign xor_ln28_63_fu_10032_p2 = (a1_192_fu_10024_p3 ^ a0_226_fu_10020_p1);

assign xor_ln28_64_fu_10046_p2 = (tmp_61_fu_10038_p3 ^ a0_225_fu_10006_p2);

assign xor_ln28_65_fu_10357_p2 = (z2_109_fu_10332_p2 ^ z1_110_fu_10326_p2);

assign xor_ln28_66_fu_10645_p2 = (z2_113_fu_10620_p2 ^ z1_114_fu_10614_p2);

assign xor_ln28_67_fu_10889_p2 = (z2_117_fu_10864_p2 ^ z1_119_fu_10858_p2);

assign xor_ln28_68_fu_10947_p2 = (a1_219_fu_10939_p3 ^ a0_244_fu_10935_p1);

assign xor_ln28_69_fu_10961_p2 = (tmp_66_fu_10953_p3 ^ a0_243_fu_10921_p2);

assign xor_ln28_6_fu_1482_p2 = (z2_10_fu_1456_p2 ^ z1_12_fu_1450_p2);

assign xor_ln28_70_fu_11195_p2 = (z2_122_fu_11170_p2 ^ z1_124_fu_11165_p2);

assign xor_ln28_71_fu_11468_p2 = (z2_126_fu_11443_p2 ^ z1_128_fu_11437_p2);

assign xor_ln28_72_fu_11760_p2 = (a1_236_fu_11752_p3 ^ a0_262_fu_11748_p1);

assign xor_ln28_73_fu_11774_p2 = (tmp_71_fu_11766_p3 ^ a0_261_fu_11734_p2);

assign xor_ln28_74_fu_11850_p2 = (a1_239_fu_11842_p3 ^ a0_265_fu_11834_p3);

assign xor_ln28_75_fu_11864_p2 = (tmp_73_fu_11856_p3 ^ a0_264_fu_11820_p1);

assign xor_ln28_76_fu_11878_p2 = (tmp_74_fu_11870_p3 ^ a0_263_fu_11806_p2);

assign xor_ln28_77_fu_12021_p2 = (z2_136_fu_11996_p2 ^ z1_137_fu_11991_p2);

assign xor_ln28_78_fu_12172_p2 = (z2_140_fu_12147_p2 ^ z1_141_fu_12142_p2);

assign xor_ln28_79_fu_12323_p2 = (z2_144_fu_12298_p2 ^ z1_146_fu_12293_p2);

assign xor_ln28_7_fu_1540_p2 = (a1_27_fu_1532_p3 ^ a0_25_fu_1528_p1);

assign xor_ln28_80_fu_12381_p2 = (a1_244_fu_12373_p3 ^ a0_270_fu_12369_p1);

assign xor_ln28_81_fu_12395_p2 = (tmp_79_fu_12387_p3 ^ a0_269_fu_12355_p2);

assign xor_ln28_82_fu_12546_p2 = (z2_149_fu_12521_p2 ^ z1_150_fu_12516_p2);

assign xor_ln28_83_fu_12697_p2 = (z2_153_fu_12672_p2 ^ z1_154_fu_12667_p2);

assign xor_ln28_84_fu_12848_p2 = (z2_157_fu_12823_p2 ^ z1_159_fu_12818_p2);

assign xor_ln28_85_fu_12906_p2 = (a1_249_fu_12898_p3 ^ a0_275_fu_12894_p1);

assign xor_ln28_86_fu_12920_p2 = (tmp_84_fu_12912_p3 ^ a0_274_fu_12880_p2);

assign xor_ln28_87_fu_13071_p2 = (z2_162_fu_13046_p2 ^ z1_164_fu_13041_p2);

assign xor_ln28_88_fu_13222_p2 = (z2_166_fu_13197_p2 ^ z1_168_fu_13192_p2);

assign xor_ln28_89_fu_13373_p2 = (z2_170_fu_13348_p2 ^ z1_173_fu_13343_p2);

assign xor_ln28_8_fu_1554_p2 = (tmp_5_fu_1546_p3 ^ a0_24_fu_1514_p2);

assign xor_ln28_90_fu_13431_p2 = (a1_254_fu_13423_p3 ^ a0_280_fu_13419_p1);

assign xor_ln28_91_fu_13445_p2 = (tmp_89_fu_13437_p3 ^ a0_279_fu_13405_p2);

assign xor_ln28_92_fu_13521_p2 = (a1_257_fu_13513_p3 ^ a0_283_fu_13505_p3);

assign xor_ln28_93_fu_13535_p2 = (tmp_91_fu_13527_p3 ^ a0_282_fu_13491_p1);

assign xor_ln28_94_fu_13549_p2 = (tmp_92_fu_13541_p3 ^ a0_281_fu_13477_p2);

assign xor_ln28_9_fu_2038_p2 = (z2_15_fu_2012_p2 ^ z1_16_fu_2006_p2);

assign xor_ln28_fu_11702_p2 = (z2_130_fu_11677_p2 ^ z1_133_fu_11672_p2);

assign xor_ln33_1_fu_5668_p2 = (trunc_ln40_1_fu_474_p4 ^ trunc_ln28_4_fu_338_p4);

assign xor_ln33_fu_1718_p2 = (xor_ln40_1_fu_490_p2 ^ trunc_ln43_1_fu_1702_p4);

assign xor_ln36_1_fu_7296_p2 = (b_185_fu_7222_p2 ^ a0_370_fu_6785_p2);

assign xor_ln36_2_fu_7302_p2 = (xor_ln45_141_fu_6962_p2 ^ a0_150_fu_7134_p2);

assign xor_ln36_fu_7290_p2 = (tmp_115_fu_7276_p3 ^ tmp_114_fu_7268_p3);

assign xor_ln40_1_fu_490_p2 = (trunc_ln70_4_fu_412_p1 ^ trunc_ln40_1_fu_474_p4);

assign xor_ln43_14_fu_1668_p2 = (trunc_ln70_4_fu_412_p1 ^ trunc_ln43_s_fu_1652_p4);

assign xor_ln43_71_fu_9227_p2 = (xor_ln45_211_fu_8719_p2 ^ a0_203_fu_8789_p2);

assign xor_ln43_83_fu_10118_p2 = (trunc_ln43_2_fu_10104_p3 ^ a0_419_cast_fu_9253_p3);

assign xor_ln43_fu_9221_p2 = (xor_ln45_231_fu_9021_p2 ^ a0_205_fu_9091_p2);

assign xor_ln45_102_fu_3832_p2 = (z1_38_fu_3744_p3 ^ z0_37_fu_3638_p3);

assign xor_ln45_103_fu_3838_p2 = (z2_184_fu_3810_p3 ^ tmp_15_fu_3824_p3);

assign xor_ln45_104_fu_4118_p2 = (xor_ln45_133_fu_4076_p2 ^ xor_ln45_132_fu_4054_p2);

assign xor_ln45_105_fu_4124_p2 = (z2_186_fu_3952_p3 ^ z0_13_fu_1616_p3);

assign xor_ln45_106_fu_5990_p2 = (z1_40_fu_5980_p2 ^ z0_40_fu_5968_p2);

assign xor_ln45_107_fu_5996_p2 = (z2_40_fu_5986_p2 ^ z0_40_fu_5968_p2);

assign xor_ln45_108_fu_6044_p2 = (z1_41_fu_6034_p2 ^ z0_42_fu_6018_p2);

assign xor_ln45_109_fu_6050_p2 = (z2_41_fu_6040_p2 ^ z0_42_fu_6018_p2);

assign xor_ln45_10_fu_986_p2 = (z1_4_fu_974_p2 ^ z0_5_fu_956_p2);

assign xor_ln45_112_fu_3904_p2 = (z1_35_fu_3552_p3 ^ z0_31_fu_3176_p3);

assign xor_ln45_113_fu_3910_p2 = (z2_185_fu_3856_p3 ^ tmp_17_fu_3896_p3);

assign xor_ln45_114_fu_6132_p2 = (xor_ln45_160_fu_6126_p2 ^ xor_ln45_155_fu_6120_p2);

assign xor_ln45_115_fu_6138_p2 = (z2_187_fu_6098_p3 ^ z0_41_fu_6002_p3);

assign xor_ln45_116_fu_6186_p2 = (z1_44_fu_6176_p2 ^ z0_45_fu_6160_p2);

assign xor_ln45_117_fu_6192_p2 = (z2_44_fu_6182_p2 ^ z0_45_fu_6160_p2);

assign xor_ln45_118_fu_6242_p2 = (z1_45_fu_6232_p2 ^ z0_47_fu_6216_p2);

assign xor_ln45_119_fu_6248_p2 = (z2_45_fu_6238_p2 ^ z0_47_fu_6216_p2);

assign xor_ln45_11_fu_992_p2 = (z2_4_fu_980_p2 ^ z0_5_fu_956_p2);

assign xor_ln45_120_fu_3916_p2 = (xor_ln45_87_fu_3546_p2 ^ xor_ln45_77_fu_3170_p2);

assign xor_ln45_121_fu_3922_p2 = (a1_304_fu_3844_p2 ^ a0_70_fu_3850_p2);

assign xor_ln45_124_fu_6330_p2 = (xor_ln45_164_fu_6324_p2 ^ xor_ln45_163_fu_6318_p2);

assign xor_ln45_125_fu_6336_p2 = (z2_188_fu_6296_p3 ^ z0_46_fu_6198_p3);

assign xor_ln45_126_fu_6372_p2 = (z1_49_fu_6362_p2 ^ z0_49_fu_6350_p2);

assign xor_ln45_127_fu_6378_p2 = (z2_48_fu_6368_p2 ^ z0_49_fu_6350_p2);

assign xor_ln45_128_fu_6426_p2 = (z1_50_fu_6416_p2 ^ z0_51_fu_6400_p2);

assign xor_ln45_129_fu_6432_p2 = (z2_49_fu_6422_p2 ^ z0_51_fu_6400_p2);

assign xor_ln45_12_fu_1092_p2 = (z1_5_fu_1080_p2 ^ z0_7_fu_1062_p2);

assign xor_ln45_130_fu_3940_p2 = (xor_ln45_121_fu_3922_p2 ^ xor_ln45_120_fu_3916_p2);

assign xor_ln45_131_fu_3946_p2 = (xor_ln45_77_fu_3170_p2 ^ a0_70_fu_3850_p2);

assign xor_ln45_132_fu_4054_p2 = (z1_26_fu_2852_p3 ^ z0_13_fu_1616_p3);

assign xor_ln45_133_fu_4076_p2 = (z2_186_fu_3952_p3 ^ tmp_20_fu_4030_p3);

assign xor_ln45_134_fu_4082_p2 = (xor_ln45_67_fu_2834_p2 ^ xor_ln45_33_fu_1598_p2);

assign xor_ln45_135_fu_4088_p2 = (a1_305_fu_3928_p2 ^ a0_73_fu_3934_p2);

assign xor_ln45_136_fu_4094_p2 = (xor_ln45_84_fu_2840_p2 ^ xor_ln45_41_fu_1610_p2);

assign xor_ln45_137_fu_4100_p2 = (xor_ln45_131_fu_3946_p2 ^ a0_74_fu_3960_p1);

assign xor_ln45_138_fu_6598_p2 = (xor_ln45_180_fu_6580_p2 ^ xor_ln45_175_fu_6574_p2);

assign xor_ln45_139_fu_6604_p2 = (z2_190_fu_6526_p3 ^ z0_44_fu_6144_p3);

assign xor_ln45_13_fu_1098_p2 = (z2_5_fu_1086_p2 ^ z0_7_fu_1062_p2);

assign xor_ln45_140_fu_6956_p2 = (z1_53_fu_6944_p2 ^ z0_53_fu_6926_p2);

assign xor_ln45_141_fu_6962_p2 = (z2_53_fu_6950_p2 ^ z0_53_fu_6926_p2);

assign xor_ln45_142_fu_7062_p2 = (z1_54_fu_7050_p2 ^ z0_55_fu_7032_p2);

assign xor_ln45_143_fu_7068_p2 = (z2_54_fu_7056_p2 ^ z0_55_fu_7032_p2);

assign xor_ln45_144_fu_4106_p2 = (tmp_99_fu_4038_p3 ^ tmp_100_fu_4046_p3);

assign xor_ln45_145_fu_4112_p2 = (tmp_102_fu_4068_p3 ^ tmp_101_fu_4060_p3);

assign xor_ln45_146_fu_4130_p2 = (xor_ln45_145_fu_4112_p2 ^ xor_ln45_144_fu_4106_p2);

assign xor_ln45_147_fu_4136_p2 = (xor_ln45_137_fu_4100_p2 ^ xor_ln45_136_fu_4094_p2);

assign xor_ln45_148_fu_7180_p2 = (xor_ln45_193_fu_7168_p2 ^ xor_ln45_192_fu_7162_p2);

assign xor_ln45_149_fu_7186_p2 = (z2_191_fu_7140_p3 ^ z0_54_fu_6968_p3);

assign xor_ln45_150_fu_7408_p2 = (z1_57_fu_7396_p2 ^ z0_57_fu_7378_p2);

assign xor_ln45_151_fu_7414_p2 = (z2_57_fu_7402_p2 ^ z0_57_fu_7378_p2);

assign xor_ln45_152_fu_4142_p2 = (xor_ln45_135_fu_4088_p2 ^ xor_ln45_134_fu_4082_p2);

assign xor_ln45_155_fu_6120_p2 = (z1_42_fu_6056_p3 ^ z0_41_fu_6002_p3);

assign xor_ln45_156_fu_7602_p2 = (z1_60_fu_7594_p2 ^ z0_60_fu_7590_p2);

assign xor_ln45_157_fu_7608_p2 = (z2_60_fu_7598_p2 ^ z0_60_fu_7590_p2);

assign xor_ln45_158_fu_7672_p2 = (z1_61_fu_7661_p2 ^ z0_62_fu_7644_p2);

assign xor_ln45_159_fu_7678_p2 = (z2_61_fu_7667_p2 ^ z0_62_fu_7644_p2);

assign xor_ln45_160_fu_6126_p2 = (z2_187_fu_6098_p3 ^ tmp_30_fu_6112_p3);

assign xor_ln45_163_fu_6318_p2 = (z1_46_fu_6254_p3 ^ z0_46_fu_6198_p3);

assign xor_ln45_164_fu_6324_p2 = (z2_188_fu_6296_p3 ^ tmp_31_fu_6310_p3);

assign xor_ln45_166_fu_7774_p2 = (z1_64_fu_7766_p2 ^ z0_64_fu_7762_p2);

assign xor_ln45_167_fu_7780_p2 = (z2_64_fu_7770_p2 ^ z0_64_fu_7762_p2);

assign xor_ln45_168_fu_7809_p2 = (z1_65_fu_7799_p2 ^ z0_66_fu_7794_p2);

assign xor_ln45_169_fu_7815_p2 = (z2_65_fu_7804_p2 ^ z0_66_fu_7794_p2);

assign xor_ln45_16_fu_1192_p2 = (z1_6_fu_1104_p3 ^ z0_6_fu_998_p3);

assign xor_ln45_171_fu_6502_p2 = (z1_51_fu_6438_p3 ^ z0_50_fu_6384_p3);

assign xor_ln45_172_fu_6508_p2 = (z2_189_fu_6480_p3 ^ tmp_32_fu_6494_p3);

assign xor_ln45_175_fu_6574_p2 = (z1_48_fu_6342_p3 ^ z0_44_fu_6144_p3);

assign xor_ln45_176_fu_7944_p2 = (z1_68_fu_7934_p2 ^ z0_68_fu_7923_p2);

assign xor_ln45_177_fu_7950_p2 = (z2_68_fu_7939_p2 ^ z0_68_fu_7923_p2);

assign xor_ln45_178_fu_8014_p2 = (z1_69_fu_8003_p2 ^ z0_70_fu_7986_p2);

assign xor_ln45_179_fu_8020_p2 = (z2_69_fu_8009_p2 ^ z0_70_fu_7986_p2);

assign xor_ln45_17_fu_1198_p2 = (z2_175_fu_1170_p3 ^ tmp_s_fu_1184_p3);

assign xor_ln45_180_fu_6580_p2 = (z2_190_fu_6526_p3 ^ tmp_34_fu_6566_p3);

assign xor_ln45_181_fu_6586_p2 = (xor_ln45_125_fu_6336_p2 ^ xor_ln45_115_fu_6138_p2);

assign xor_ln45_182_fu_6592_p2 = (a1_332_fu_6514_p2 ^ a0_129_fu_6520_p2);

assign xor_ln45_183_fu_6610_p2 = (xor_ln45_182_fu_6592_p2 ^ xor_ln45_181_fu_6586_p2);

assign xor_ln45_184_fu_8109_p2 = (xor_ln45_236_fu_8103_p2 ^ xor_ln45_235_fu_8097_p2);

assign xor_ln45_185_fu_8115_p2 = (z2_194_fu_8075_p3 ^ z0_69_fu_7956_p3);

assign xor_ln45_186_fu_8201_p2 = (z1_72_fu_8190_p2 ^ z0_73_fu_8173_p2);

assign xor_ln45_187_fu_8207_p2 = (z2_72_fu_8196_p2 ^ z0_73_fu_8173_p2);

assign xor_ln45_188_fu_8282_p2 = (z1_73_fu_8271_p2 ^ z0_75_fu_8254_p2);

assign xor_ln45_189_fu_8288_p2 = (z2_73_fu_8277_p2 ^ z0_75_fu_8254_p2);

assign xor_ln45_18_fu_1204_p2 = (xor_ln45_17_fu_1198_p2 ^ xor_ln45_16_fu_1192_p2);

assign xor_ln45_192_fu_7162_p2 = (z1_55_fu_7074_p3 ^ z0_54_fu_6968_p3);

assign xor_ln45_193_fu_7168_p2 = (z2_191_fu_7140_p3 ^ tmp_40_fu_7154_p3);

assign xor_ln45_194_fu_8382_p2 = (xor_ln45_240_fu_8376_p2 ^ xor_ln45_239_fu_8370_p2);

assign xor_ln45_195_fu_8388_p2 = (z2_195_fu_8348_p3 ^ z0_74_fu_8213_p3);

assign xor_ln45_196_fu_8431_p2 = (z1_77_fu_8421_p2 ^ z0_77_fu_8410_p2);

assign xor_ln45_197_fu_8437_p2 = (z2_76_fu_8426_p2 ^ z0_77_fu_8410_p2);

assign xor_ln45_198_fu_8507_p2 = (z1_78_fu_8496_p2 ^ z0_79_fu_8479_p2);

assign xor_ln45_199_fu_8513_p2 = (z2_77_fu_8502_p2 ^ z0_79_fu_8479_p2);

assign xor_ln45_19_fu_1210_p2 = (z2_175_fu_1170_p3 ^ z0_6_fu_998_p3);

assign xor_ln45_1_fu_616_p2 = (z2_fu_604_p2 ^ z0_fu_580_p2);

assign xor_ln45_200_fu_7174_p2 = (xor_ln45_143_fu_7068_p2 ^ xor_ln45_141_fu_6962_p2);

assign xor_ln45_201_fu_7192_p2 = (xor_ln45_200_fu_7174_p2 ^ xor_ln28_46_fu_7148_p2);

assign xor_ln45_208_fu_7738_p2 = (z1_62_fu_7684_p3 ^ z0_61_fu_7614_p3);

assign xor_ln45_209_fu_7744_p2 = (z2_192_fu_7716_p3 ^ tmp_46_fu_7730_p3);

assign xor_ln45_20_fu_1290_p2 = (z1_9_fu_1278_p2 ^ z0_9_fu_1260_p2);

assign xor_ln45_210_fu_8713_p2 = (z1_81_fu_8703_p2 ^ z0_81_fu_8698_p2);

assign xor_ln45_211_fu_8719_p2 = (z2_81_fu_8708_p2 ^ z0_81_fu_8698_p2);

assign xor_ln45_212_fu_8748_p2 = (z1_82_fu_8738_p2 ^ z0_83_fu_8733_p2);

assign xor_ln45_213_fu_8754_p2 = (z2_82_fu_8743_p2 ^ z0_83_fu_8733_p2);

assign xor_ln45_218_fu_8829_p2 = (xor_ln45_272_fu_8823_p2 ^ xor_ln45_271_fu_8817_p2);

assign xor_ln45_219_fu_8835_p2 = (z2_198_fu_8795_p3 ^ z0_82_fu_8725_p3);

assign xor_ln45_21_fu_1296_p2 = (z2_8_fu_1284_p2 ^ z0_9_fu_1260_p2);

assign xor_ln45_220_fu_8864_p2 = (z1_85_fu_8854_p2 ^ z0_86_fu_8849_p2);

assign xor_ln45_221_fu_8870_p2 = (z2_85_fu_8859_p2 ^ z0_86_fu_8849_p2);

assign xor_ln45_222_fu_8899_p2 = (z1_86_fu_8889_p2 ^ z0_88_fu_8884_p2);

assign xor_ln45_223_fu_8905_p2 = (z2_86_fu_8894_p2 ^ z0_88_fu_8884_p2);

assign xor_ln45_228_fu_8980_p2 = (xor_ln45_282_fu_8974_p2 ^ xor_ln45_275_fu_8968_p2);

assign xor_ln45_229_fu_8986_p2 = (z2_199_fu_8946_p3 ^ z0_87_fu_8876_p3);

assign xor_ln45_22_fu_1396_p2 = (z1_10_fu_1384_p2 ^ z0_11_fu_1366_p2);

assign xor_ln45_230_fu_9015_p2 = (z1_90_fu_9005_p2 ^ z0_90_fu_9000_p2);

assign xor_ln45_231_fu_9021_p2 = (z2_89_fu_9010_p2 ^ z0_90_fu_9000_p2);

assign xor_ln45_232_fu_9050_p2 = (z1_91_fu_9040_p2 ^ z0_92_fu_9035_p2);

assign xor_ln45_233_fu_9056_p2 = (z2_90_fu_9045_p2 ^ z0_92_fu_9035_p2);

assign xor_ln45_235_fu_8097_p2 = (z1_70_fu_8026_p3 ^ z0_69_fu_7956_p3);

assign xor_ln45_236_fu_8103_p2 = (z2_194_fu_8075_p3 ^ tmp_48_fu_8089_p3);

assign xor_ln45_239_fu_8370_p2 = (z1_74_fu_8294_p3 ^ z0_74_fu_8213_p3);

assign xor_ln45_23_fu_1402_p2 = (z2_9_fu_1390_p2 ^ z0_11_fu_1366_p2);

assign xor_ln45_240_fu_8376_p2 = (z2_195_fu_8348_p3 ^ tmp_49_fu_8362_p3);

assign xor_ln45_243_fu_8590_p2 = (z1_79_fu_8519_p3 ^ z0_78_fu_8443_p3);

assign xor_ln45_244_fu_9320_p2 = (z1_94_fu_9310_p2 ^ z0_94_fu_9299_p2);

assign xor_ln45_245_fu_9326_p2 = (z2_94_fu_9315_p2 ^ z0_94_fu_9299_p2);

assign xor_ln45_246_fu_9400_p2 = (z1_95_fu_9389_p2 ^ z0_96_fu_9372_p2);

assign xor_ln45_247_fu_9406_p2 = (z2_95_fu_9395_p2 ^ z0_96_fu_9372_p2);

assign xor_ln45_248_fu_8596_p2 = (z2_196_fu_8568_p3 ^ tmp_50_fu_8582_p3);

assign xor_ln45_251_fu_8662_p2 = (z1_76_fu_8394_p3 ^ z0_72_fu_8121_p3);

assign xor_ln45_252_fu_9495_p2 = (xor_ln45_316_fu_9489_p2 ^ xor_ln45_309_fu_9483_p2);

assign xor_ln45_253_fu_9501_p2 = (z2_202_fu_9461_p3 ^ z0_95_fu_9332_p3);

assign xor_ln45_254_fu_9585_p2 = (z1_98_fu_9574_p2 ^ z0_99_fu_9557_p2);

assign xor_ln45_255_fu_9591_p2 = (z2_98_fu_9580_p2 ^ z0_99_fu_9557_p2);

assign xor_ln45_256_fu_9666_p2 = (z1_99_fu_9655_p2 ^ z0_101_fu_9638_p2);

assign xor_ln45_257_fu_9672_p2 = (z2_99_fu_9661_p2 ^ z0_101_fu_9638_p2);

assign xor_ln45_258_fu_8668_p2 = (z2_197_fu_8614_p3 ^ tmp_52_fu_8654_p3);

assign xor_ln45_259_fu_8674_p2 = (xor_ln45_195_fu_8388_p2 ^ xor_ln45_185_fu_8115_p2);

assign xor_ln45_260_fu_8680_p2 = (a1_364_fu_8602_p2 ^ a0_201_fu_8608_p2);

assign xor_ln45_262_fu_9766_p2 = (xor_ln45_326_fu_9760_p2 ^ xor_ln45_319_fu_9754_p2);

assign xor_ln45_263_fu_9772_p2 = (z2_203_fu_9732_p3 ^ z0_100_fu_9597_p3);

assign xor_ln45_264_fu_9825_p2 = (z1_103_fu_9815_p2 ^ z0_103_fu_9804_p2);

assign xor_ln45_265_fu_9831_p2 = (z2_102_fu_9820_p2 ^ z0_103_fu_9804_p2);

assign xor_ln45_266_fu_9905_p2 = (z1_104_fu_9894_p2 ^ z0_105_fu_9877_p2);

assign xor_ln45_267_fu_9911_p2 = (z2_103_fu_9900_p2 ^ z0_105_fu_9877_p2);

assign xor_ln45_26_fu_1496_p2 = (z1_11_fu_1408_p3 ^ z0_10_fu_1302_p3);

assign xor_ln45_271_fu_8817_p2 = (z1_83_fu_8760_p3 ^ z0_82_fu_8725_p3);

assign xor_ln45_272_fu_8823_p2 = (z2_198_fu_8795_p3 ^ tmp_53_fu_8809_p3);

assign xor_ln45_275_fu_8968_p2 = (z1_87_fu_8911_p3 ^ z0_87_fu_8876_p3);

assign xor_ln45_276_fu_10072_p2 = (xor_ln45_340_fu_10066_p2 ^ xor_ln45_339_fu_10060_p2);

assign xor_ln45_277_fu_10078_p2 = (z2_205_fu_10012_p3 ^ z0_98_fu_9507_p3);

assign xor_ln45_278_fu_10202_p2 = (z1_107_fu_10191_p2 ^ z0_108_fu_10174_p2);

assign xor_ln45_279_fu_10208_p2 = (z2_107_fu_10197_p2 ^ z0_108_fu_10174_p2);

assign xor_ln45_27_fu_1502_p2 = (z2_176_fu_1474_p3 ^ tmp_4_fu_1488_p3);

assign xor_ln45_280_fu_10283_p2 = (z1_108_fu_10272_p2 ^ z0_110_fu_10255_p2);

assign xor_ln45_281_fu_10289_p2 = (z2_108_fu_10278_p2 ^ z0_110_fu_10255_p2);

assign xor_ln45_282_fu_8974_p2 = (z2_199_fu_8946_p3 ^ tmp_54_fu_8960_p3);

assign xor_ln45_285_fu_9119_p2 = (z1_92_fu_9062_p3 ^ z0_91_fu_9027_p3);

assign xor_ln45_286_fu_10383_p2 = (xor_ln45_344_fu_10377_p2 ^ xor_ln45_343_fu_10371_p2);

assign xor_ln45_287_fu_10389_p2 = (z2_206_fu_10349_p3 ^ z0_109_fu_10214_p3);

assign xor_ln45_288_fu_10490_p2 = (z1_111_fu_10479_p2 ^ z0_113_fu_10462_p2);

assign xor_ln45_289_fu_10496_p2 = (z2_111_fu_10485_p2 ^ z0_113_fu_10462_p2);

assign xor_ln45_290_fu_10571_p2 = (z1_112_fu_10560_p2 ^ z0_115_fu_10543_p2);

assign xor_ln45_291_fu_10577_p2 = (z2_112_fu_10566_p2 ^ z0_115_fu_10543_p2);

assign xor_ln45_292_fu_9125_p2 = (z2_200_fu_9097_p3 ^ tmp_55_fu_9111_p3);

assign xor_ln45_296_fu_10671_p2 = (xor_ln45_354_fu_10665_p2 ^ xor_ln45_347_fu_10659_p2);

assign xor_ln45_297_fu_10677_p2 = (z2_207_fu_10637_p3 ^ z0_114_fu_10502_p3);

assign xor_ln45_298_fu_10735_p2 = (z1_116_fu_10724_p2 ^ z0_117_fu_10709_p2);

assign xor_ln45_299_fu_10741_p2 = (z2_115_fu_10730_p2 ^ z0_117_fu_10709_p2);

assign xor_ln45_2_fu_716_p2 = (z1_1_fu_704_p2 ^ z0_2_fu_686_p2);

assign xor_ln45_300_fu_10815_p2 = (z1_117_fu_10804_p2 ^ z0_119_fu_10787_p2);

assign xor_ln45_301_fu_10821_p2 = (z2_116_fu_10810_p2 ^ z0_119_fu_10787_p2);

assign xor_ln45_304_fu_9209_p2 = (xor_ln45_229_fu_8986_p2 ^ a1_365_fu_9131_p2);

assign xor_ln45_306_fu_9239_p2 = (xor_ln45_304_fu_9209_p2 ^ a0_395_fu_9203_p2);

assign xor_ln45_309_fu_9483_p2 = (z1_96_fu_9412_p3 ^ z0_95_fu_9332_p3);

assign xor_ln45_30_fu_1568_p2 = (z1_8_fu_1216_p3 ^ z0_4_fu_840_p3);

assign xor_ln45_310_fu_10987_p2 = (xor_ln45_374_fu_10981_p2 ^ xor_ln45_367_fu_10975_p2);

assign xor_ln45_311_fu_10993_p2 = (z2_209_fu_10927_p3 ^ z0_112_fu_10395_p3);

assign xor_ln45_312_fu_11046_p2 = (z1_121_fu_11036_p2 ^ z0_121_fu_11025_p2);

assign xor_ln45_313_fu_11052_p2 = (z2_120_fu_11041_p2 ^ z0_121_fu_11025_p2);

assign xor_ln45_314_fu_11126_p2 = (z1_122_fu_11115_p2 ^ z0_123_fu_11098_p2);

assign xor_ln45_315_fu_11132_p2 = (z2_121_fu_11121_p2 ^ z0_123_fu_11098_p2);

assign xor_ln45_316_fu_9489_p2 = (z2_202_fu_9461_p3 ^ tmp_58_fu_9475_p3);

assign xor_ln45_319_fu_9754_p2 = (z1_100_fu_9678_p3 ^ z0_100_fu_9597_p3);

assign xor_ln45_31_fu_1574_p2 = (z2_177_fu_1520_p3 ^ tmp_6_fu_1560_p3);

assign xor_ln45_320_fu_11221_p2 = (xor_ln45_378_fu_11215_p2 ^ xor_ln45_377_fu_11209_p2);

assign xor_ln45_321_fu_11227_p2 = (z2_210_fu_11187_p3 ^ z0_122_fu_11058_p3);

assign xor_ln45_322_fu_11313_p2 = (z1_125_fu_11302_p2 ^ z0_126_fu_11285_p2);

assign xor_ln45_323_fu_11319_p2 = (z2_124_fu_11308_p2 ^ z0_126_fu_11285_p2);

assign xor_ln45_324_fu_11394_p2 = (z1_126_fu_11383_p2 ^ z0_128_fu_11366_p2);

assign xor_ln45_325_fu_11400_p2 = (z2_125_fu_11389_p2 ^ z0_128_fu_11366_p2);

assign xor_ln45_326_fu_9760_p2 = (z2_203_fu_9732_p3 ^ tmp_59_fu_9746_p3);

assign xor_ln45_329_fu_9988_p2 = (z1_105_fu_9917_p3 ^ z0_104_fu_9837_p3);

assign xor_ln45_32_fu_1592_p2 = (xor_ln45_31_fu_1574_p2 ^ xor_ln45_30_fu_1568_p2);

assign xor_ln45_330_fu_11494_p2 = (xor_ln45_388_fu_11488_p2 ^ xor_ln45_381_fu_11482_p2);

assign xor_ln45_331_fu_11500_p2 = (z2_211_fu_11460_p3 ^ z0_127_fu_11325_p3);

assign xor_ln45_332_fu_11553_p2 = (z1_130_fu_11543_p2 ^ z0_130_fu_11532_p2);

assign xor_ln45_333_fu_11559_p2 = (z2_128_fu_11548_p2 ^ z0_130_fu_11532_p2);

assign xor_ln45_334_fu_11633_p2 = (z1_131_fu_11622_p2 ^ z0_132_fu_11605_p2);

assign xor_ln45_335_fu_11639_p2 = (z2_129_fu_11628_p2 ^ z0_132_fu_11605_p2);

assign xor_ln45_336_fu_9994_p2 = (z2_204_fu_9966_p3 ^ tmp_60_fu_9980_p3);

assign xor_ln45_339_fu_10060_p2 = (z1_102_fu_9778_p3 ^ z0_98_fu_9507_p3);

assign xor_ln45_33_fu_1598_p2 = (z2_177_fu_1520_p3 ^ z0_4_fu_840_p3);

assign xor_ln45_340_fu_10066_p2 = (z2_205_fu_10012_p3 ^ tmp_62_fu_10052_p3);

assign xor_ln45_343_fu_10371_p2 = (z1_109_fu_10295_p3 ^ z0_109_fu_10214_p3);

assign xor_ln45_344_fu_10377_p2 = (z2_206_fu_10349_p3 ^ tmp_63_fu_10363_p3);

assign xor_ln45_347_fu_10659_p2 = (z1_113_fu_10583_p3 ^ z0_114_fu_10502_p3);

assign xor_ln45_348_fu_11904_p2 = (xor_ln45_412_fu_11898_p2 ^ xor_ln45_411_fu_11892_p2);

assign xor_ln45_349_fu_11910_p2 = (z2_214_fu_11812_p3 ^ z0_107_fu_10084_p3);

assign xor_ln45_34_fu_1846_p2 = (z1_13_fu_1834_p2 ^ z0_14_fu_1816_p2);

assign xor_ln45_350_fu_11931_p2 = (z1_134_fu_11921_p2 ^ z0_134_fu_11916_p2);

assign xor_ln45_351_fu_11937_p2 = (z2_134_fu_11926_p2 ^ z0_134_fu_11916_p2);

assign xor_ln45_352_fu_11966_p2 = (z1_135_fu_11956_p2 ^ z0_136_fu_11951_p2);

assign xor_ln45_353_fu_11972_p2 = (z2_135_fu_11961_p2 ^ z0_136_fu_11951_p2);

assign xor_ln45_354_fu_10665_p2 = (z2_207_fu_10637_p3 ^ tmp_64_fu_10651_p3);

assign xor_ln45_357_fu_10903_p2 = (z1_118_fu_10827_p3 ^ z0_118_fu_10747_p3);

assign xor_ln45_358_fu_12047_p2 = (xor_ln45_422_fu_12041_p2 ^ xor_ln45_415_fu_12035_p2);

assign xor_ln45_359_fu_12053_p2 = (z2_215_fu_12013_p3 ^ z0_135_fu_11943_p3);

assign xor_ln45_35_fu_1852_p2 = (z2_13_fu_1840_p2 ^ z0_14_fu_1816_p2);

assign xor_ln45_360_fu_12082_p2 = (z1_138_fu_12072_p2 ^ z0_139_fu_12067_p2);

assign xor_ln45_361_fu_12088_p2 = (z2_138_fu_12077_p2 ^ z0_139_fu_12067_p2);

assign xor_ln45_362_fu_12117_p2 = (z1_139_fu_12107_p2 ^ z0_141_fu_12102_p2);

assign xor_ln45_363_fu_12123_p2 = (z2_139_fu_12112_p2 ^ z0_141_fu_12102_p2);

assign xor_ln45_364_fu_10909_p2 = (z2_208_fu_10881_p3 ^ tmp_65_fu_10895_p3);

assign xor_ln45_367_fu_10975_p2 = (z1_115_fu_10683_p3 ^ z0_112_fu_10395_p3);

assign xor_ln45_368_fu_12198_p2 = (xor_ln45_432_fu_12192_p2 ^ xor_ln45_425_fu_12186_p2);

assign xor_ln45_369_fu_12204_p2 = (z2_216_fu_12164_p3 ^ z0_140_fu_12094_p3);

assign xor_ln45_36_fu_1952_p2 = (z1_14_fu_1940_p2 ^ z0_16_fu_1922_p2);

assign xor_ln45_370_fu_12233_p2 = (z1_143_fu_12223_p2 ^ z0_143_fu_12218_p2);

assign xor_ln45_371_fu_12239_p2 = (z2_142_fu_12228_p2 ^ z0_143_fu_12218_p2);

assign xor_ln45_372_fu_12268_p2 = (z1_144_fu_12258_p2 ^ z0_145_fu_12253_p2);

assign xor_ln45_373_fu_12274_p2 = (z2_143_fu_12263_p2 ^ z0_145_fu_12253_p2);

assign xor_ln45_374_fu_10981_p2 = (z2_209_fu_10927_p3 ^ tmp_67_fu_10967_p3);

assign xor_ln45_377_fu_11209_p2 = (z1_123_fu_11138_p3 ^ z0_122_fu_11058_p3);

assign xor_ln45_378_fu_11215_p2 = (z2_210_fu_11187_p3 ^ tmp_68_fu_11201_p3);

assign xor_ln45_37_fu_1958_p2 = (z2_14_fu_1946_p2 ^ z0_16_fu_1922_p2);

assign xor_ln45_381_fu_11482_p2 = (z1_127_fu_11406_p3 ^ z0_127_fu_11325_p3);

assign xor_ln45_382_fu_12421_p2 = (xor_ln45_446_fu_12415_p2 ^ xor_ln45_445_fu_12409_p2);

assign xor_ln45_383_fu_12427_p2 = (z2_218_fu_12361_p3 ^ z0_138_fu_12059_p3);

assign xor_ln45_384_fu_12456_p2 = (z1_147_fu_12446_p2 ^ z0_148_fu_12441_p2);

assign xor_ln45_385_fu_12462_p2 = (z2_147_fu_12451_p2 ^ z0_148_fu_12441_p2);

assign xor_ln45_386_fu_12491_p2 = (z1_148_fu_12481_p2 ^ z0_150_fu_12476_p2);

assign xor_ln45_387_fu_12497_p2 = (z2_148_fu_12486_p2 ^ z0_150_fu_12476_p2);

assign xor_ln45_388_fu_11488_p2 = (z2_211_fu_11460_p3 ^ tmp_69_fu_11474_p3);

assign xor_ln45_38_fu_1580_p2 = (xor_ln45_9_fu_834_p2 ^ xor_ln45_19_fu_1210_p2);

assign xor_ln45_391_fu_11716_p2 = (z1_132_fu_11645_p3 ^ z0_131_fu_11565_p3);

assign xor_ln45_392_fu_12572_p2 = (xor_ln45_450_fu_12566_p2 ^ xor_ln45_449_fu_12560_p2);

assign xor_ln45_393_fu_12578_p2 = (z2_219_fu_12538_p3 ^ z0_149_fu_12468_p3);

assign xor_ln45_394_fu_12607_p2 = (z1_151_fu_12597_p2 ^ z0_153_fu_12592_p2);

assign xor_ln45_395_fu_12613_p2 = (z2_151_fu_12602_p2 ^ z0_153_fu_12592_p2);

assign xor_ln45_396_fu_12642_p2 = (z1_152_fu_12632_p2 ^ z0_155_fu_12627_p2);

assign xor_ln45_397_fu_12648_p2 = (z2_152_fu_12637_p2 ^ z0_155_fu_12627_p2);

assign xor_ln45_398_fu_11722_p2 = (z2_212_fu_11694_p3 ^ tmp_70_fu_11708_p3);

assign xor_ln45_39_fu_1586_p2 = (a1_276_fu_1508_p2 ^ a0_24_fu_1514_p2);

assign xor_ln45_3_fu_722_p2 = (z2_1_fu_710_p2 ^ z0_2_fu_686_p2);

assign xor_ln45_401_fu_11788_p2 = (z1_129_fu_11506_p3 ^ z0_125_fu_11233_p3);

assign xor_ln45_402_fu_12723_p2 = (xor_ln45_456_fu_12717_p2 ^ xor_ln45_453_fu_12711_p2);

assign xor_ln45_403_fu_12729_p2 = (z2_220_fu_12689_p3 ^ z0_154_fu_12619_p3);

assign xor_ln45_404_fu_12758_p2 = (z1_156_fu_12748_p2 ^ z0_157_fu_12743_p2);

assign xor_ln45_405_fu_12764_p2 = (z2_155_fu_12753_p2 ^ z0_157_fu_12743_p2);

assign xor_ln45_406_fu_12793_p2 = (z1_157_fu_12783_p2 ^ z0_159_fu_12778_p2);

assign xor_ln45_407_fu_12799_p2 = (z2_156_fu_12788_p2 ^ z0_159_fu_12778_p2);

assign xor_ln45_408_fu_11794_p2 = (z2_213_fu_11740_p3 ^ tmp_72_fu_11780_p3);

assign xor_ln45_40_fu_1604_p2 = (xor_ln45_39_fu_1586_p2 ^ xor_ln45_38_fu_1580_p2);

assign xor_ln45_411_fu_11892_p2 = (z1_120_fu_10999_p3 ^ z0_107_fu_10084_p3);

assign xor_ln45_412_fu_11898_p2 = (z2_214_fu_11812_p3 ^ tmp_75_fu_11884_p3);

assign xor_ln45_415_fu_12035_p2 = (z1_136_fu_11978_p3 ^ z0_135_fu_11943_p3);

assign xor_ln45_416_fu_12946_p2 = (xor_ln45_464_fu_12940_p2 ^ xor_ln45_463_fu_12934_p2);

assign xor_ln45_417_fu_12952_p2 = (z2_222_fu_12886_p3 ^ z0_152_fu_12584_p3);

assign xor_ln45_418_fu_12981_p2 = (z1_161_fu_12971_p2 ^ z0_161_fu_12966_p2);

assign xor_ln45_419_fu_12987_p2 = (z2_160_fu_12976_p2 ^ z0_161_fu_12966_p2);

assign xor_ln45_41_fu_1610_p2 = (xor_ln45_9_fu_834_p2 ^ a0_24_fu_1514_p2);

assign xor_ln45_420_fu_13016_p2 = (z1_162_fu_13006_p2 ^ z0_163_fu_13001_p2);

assign xor_ln45_421_fu_13022_p2 = (z2_161_fu_13011_p2 ^ z0_163_fu_13001_p2);

assign xor_ln45_422_fu_12041_p2 = (z2_215_fu_12013_p3 ^ tmp_76_fu_12027_p3);

assign xor_ln45_425_fu_12186_p2 = (z1_140_fu_12129_p3 ^ z0_140_fu_12094_p3);

assign xor_ln45_426_fu_13097_p2 = (xor_ln45_468_fu_13091_p2 ^ xor_ln45_467_fu_13085_p2);

assign xor_ln45_427_fu_13103_p2 = (z2_223_fu_13063_p3 ^ z0_162_fu_12993_p3);

assign xor_ln45_428_fu_13132_p2 = (z1_165_fu_13122_p2 ^ z0_166_fu_13117_p2);

assign xor_ln45_429_fu_13138_p2 = (z2_164_fu_13127_p2 ^ z0_166_fu_13117_p2);

assign xor_ln45_42_fu_2064_p2 = (xor_ln45_51_fu_2058_p2 ^ xor_ln45_50_fu_2052_p2);

assign xor_ln45_430_fu_13167_p2 = (z1_166_fu_13157_p2 ^ z0_168_fu_13152_p2);

assign xor_ln45_431_fu_13173_p2 = (z2_165_fu_13162_p2 ^ z0_168_fu_13152_p2);

assign xor_ln45_432_fu_12192_p2 = (z2_216_fu_12164_p3 ^ tmp_77_fu_12178_p3);

assign xor_ln45_435_fu_12337_p2 = (z1_145_fu_12280_p3 ^ z0_144_fu_12245_p3);

assign xor_ln45_436_fu_13248_p2 = (xor_ln45_472_fu_13242_p2 ^ xor_ln45_471_fu_13236_p2);

assign xor_ln45_437_fu_13254_p2 = (z2_224_fu_13214_p3 ^ z0_167_fu_13144_p3);

assign xor_ln45_438_fu_13283_p2 = (z1_170_fu_13273_p2 ^ z0_170_fu_13268_p2);

assign xor_ln45_439_fu_13289_p2 = (z2_168_fu_13278_p2 ^ z0_170_fu_13268_p2);

assign xor_ln45_43_fu_2070_p2 = (z2_178_fu_2030_p3 ^ z0_15_fu_1858_p3);

assign xor_ln45_440_fu_13318_p2 = (z1_171_fu_13308_p2 ^ z0_172_fu_13303_p2);

assign xor_ln45_441_fu_13324_p2 = (z2_169_fu_13313_p2 ^ z0_172_fu_13303_p2);

assign xor_ln45_442_fu_12343_p2 = (z2_217_fu_12315_p3 ^ tmp_78_fu_12329_p3);

assign xor_ln45_445_fu_12409_p2 = (z1_142_fu_12210_p3 ^ z0_138_fu_12059_p3);

assign xor_ln45_446_fu_12415_p2 = (z2_218_fu_12361_p3 ^ tmp_80_fu_12401_p3);

assign xor_ln45_449_fu_12560_p2 = (z1_149_fu_12503_p3 ^ z0_149_fu_12468_p3);

assign xor_ln45_44_fu_2222_p2 = (z1_17_fu_2210_p2 ^ z0_19_fu_2192_p2);

assign xor_ln45_450_fu_12566_p2 = (z2_219_fu_12538_p3 ^ tmp_81_fu_12552_p3);

assign xor_ln45_453_fu_12711_p2 = (z1_153_fu_12654_p3 ^ z0_154_fu_12619_p3);

assign xor_ln45_454_fu_13575_p2 = (xor_ln45_484_fu_13569_p2 ^ xor_ln45_483_fu_13563_p2);

assign xor_ln45_455_fu_13581_p2 = (z2_227_fu_13483_p3 ^ z0_147_fu_12433_p3);

assign xor_ln45_456_fu_12717_p2 = (z2_220_fu_12689_p3 ^ tmp_82_fu_12703_p3);

assign xor_ln45_459_fu_12862_p2 = (z1_158_fu_12805_p3 ^ z0_158_fu_12770_p3);

assign xor_ln45_45_fu_2228_p2 = (z2_17_fu_2216_p2 ^ z0_19_fu_2192_p2);

assign xor_ln45_460_fu_12868_p2 = (z2_221_fu_12840_p3 ^ tmp_83_fu_12854_p3);

assign xor_ln45_463_fu_12934_p2 = (z1_155_fu_12735_p3 ^ z0_152_fu_12584_p3);

assign xor_ln45_464_fu_12940_p2 = (z2_222_fu_12886_p3 ^ tmp_85_fu_12926_p3);

assign xor_ln45_467_fu_13085_p2 = (z1_163_fu_13028_p3 ^ z0_162_fu_12993_p3);

assign xor_ln45_468_fu_13091_p2 = (z2_223_fu_13063_p3 ^ tmp_86_fu_13077_p3);

assign xor_ln45_46_fu_2328_p2 = (z1_18_fu_2316_p2 ^ z0_21_fu_2298_p2);

assign xor_ln45_471_fu_13236_p2 = (z1_167_fu_13179_p3 ^ z0_167_fu_13144_p3);

assign xor_ln45_472_fu_13242_p2 = (z2_224_fu_13214_p3 ^ tmp_87_fu_13228_p3);

assign xor_ln45_475_fu_13387_p2 = (z1_172_fu_13330_p3 ^ z0_171_fu_13295_p3);

assign xor_ln45_476_fu_13393_p2 = (z2_225_fu_13365_p3 ^ tmp_88_fu_13379_p3);

assign xor_ln45_479_fu_13459_p2 = (z1_169_fu_13260_p3 ^ z0_165_fu_13109_p3);

assign xor_ln45_47_fu_2334_p2 = (z2_18_fu_2322_p2 ^ z0_21_fu_2298_p2);

assign xor_ln45_480_fu_13465_p2 = (z2_226_fu_13411_p3 ^ tmp_90_fu_13451_p3);

assign xor_ln45_483_fu_13563_p2 = (z1_160_fu_12958_p3 ^ z0_147_fu_12433_p3);

assign xor_ln45_484_fu_13569_p2 = (z2_227_fu_13483_p3 ^ tmp_93_fu_13555_p3);

assign xor_ln45_50_fu_2052_p2 = (z1_15_fu_1964_p3 ^ z0_15_fu_1858_p3);

assign xor_ln45_51_fu_2058_p2 = (z2_178_fu_2030_p3 ^ tmp_8_fu_2044_p3);

assign xor_ln45_52_fu_2440_p2 = (xor_ln45_61_fu_2434_p2 ^ xor_ln45_60_fu_2428_p2);

assign xor_ln45_53_fu_2446_p2 = (z2_179_fu_2406_p3 ^ z0_20_fu_2234_p3);

assign xor_ln45_54_fu_2526_p2 = (z1_22_fu_2514_p2 ^ z0_23_fu_2496_p2);

assign xor_ln45_55_fu_2532_p2 = (z2_21_fu_2520_p2 ^ z0_23_fu_2496_p2);

assign xor_ln45_56_fu_2632_p2 = (z1_23_fu_2620_p2 ^ z0_25_fu_2602_p2);

assign xor_ln45_57_fu_2638_p2 = (z2_22_fu_2626_p2 ^ z0_25_fu_2602_p2);

assign xor_ln45_60_fu_2428_p2 = (z1_19_fu_2340_p3 ^ z0_20_fu_2234_p3);

assign xor_ln45_61_fu_2434_p2 = (z2_179_fu_2406_p3 ^ tmp_9_fu_2420_p3);

assign xor_ln45_64_fu_2732_p2 = (z1_24_fu_2644_p3 ^ z0_24_fu_2538_p3);

assign xor_ln45_65_fu_2738_p2 = (z2_180_fu_2710_p3 ^ tmp_10_fu_2724_p3);

assign xor_ln45_66_fu_2828_p2 = (xor_ln45_75_fu_2810_p2 ^ xor_ln45_74_fu_2804_p2);

assign xor_ln45_67_fu_2834_p2 = (z2_181_fu_2756_p3 ^ z0_18_fu_2076_p3);

assign xor_ln45_68_fu_2946_p2 = (z1_27_fu_2934_p2 ^ z0_27_fu_2916_p2);

assign xor_ln45_69_fu_2952_p2 = (z2_26_fu_2940_p2 ^ z0_27_fu_2916_p2);

assign xor_ln45_6_fu_816_p2 = (z1_2_fu_728_p3 ^ z0_1_fu_622_p3);

assign xor_ln45_70_fu_3052_p2 = (z1_28_fu_3040_p2 ^ z0_29_fu_3022_p2);

assign xor_ln45_71_fu_3058_p2 = (z2_27_fu_3046_p2 ^ z0_29_fu_3022_p2);

assign xor_ln45_74_fu_2804_p2 = (z1_21_fu_2452_p3 ^ z0_18_fu_2076_p3);

assign xor_ln45_75_fu_2810_p2 = (z2_181_fu_2756_p3 ^ tmp_12_fu_2796_p3);

assign xor_ln45_76_fu_3164_p2 = (xor_ln45_95_fu_3158_p2 ^ xor_ln45_94_fu_3152_p2);

assign xor_ln45_77_fu_3170_p2 = (z2_182_fu_3130_p3 ^ z0_28_fu_2958_p3);

assign xor_ln45_78_fu_3322_p2 = (z1_31_fu_3310_p2 ^ z0_32_fu_3292_p2);

assign xor_ln45_79_fu_3328_p2 = (z2_30_fu_3316_p2 ^ z0_32_fu_3292_p2);

assign xor_ln45_7_fu_822_p2 = (z2_174_fu_794_p3 ^ tmp_7_fu_808_p3);

assign xor_ln45_80_fu_3428_p2 = (z1_32_fu_3416_p2 ^ z0_34_fu_3398_p2);

assign xor_ln45_81_fu_3434_p2 = (z2_31_fu_3422_p2 ^ z0_34_fu_3398_p2);

assign xor_ln45_82_fu_2816_p2 = (xor_ln45_53_fu_2446_p2 ^ xor_ln45_43_fu_2070_p2);

assign xor_ln45_83_fu_2822_p2 = (a1_290_fu_2744_p2 ^ a0_50_fu_2750_p2);

assign xor_ln45_84_fu_2840_p2 = (xor_ln45_43_fu_2070_p2 ^ a0_50_fu_2750_p2);

assign xor_ln45_85_fu_2846_p2 = (xor_ln45_83_fu_2822_p2 ^ xor_ln45_82_fu_2816_p2);

assign xor_ln45_86_fu_3540_p2 = (xor_ln45_99_fu_3534_p2 ^ xor_ln45_98_fu_3528_p2);

assign xor_ln45_87_fu_3546_p2 = (z2_183_fu_3506_p3 ^ z0_33_fu_3334_p3);

assign xor_ln45_88_fu_3626_p2 = (z1_36_fu_3614_p2 ^ z0_36_fu_3596_p2);

assign xor_ln45_89_fu_3632_p2 = (z2_34_fu_3620_p2 ^ z0_36_fu_3596_p2);

assign xor_ln45_8_fu_828_p2 = (xor_ln45_7_fu_822_p2 ^ xor_ln45_6_fu_816_p2);

assign xor_ln45_90_fu_3732_p2 = (z1_37_fu_3720_p2 ^ z0_38_fu_3702_p2);

assign xor_ln45_91_fu_3738_p2 = (z2_35_fu_3726_p2 ^ z0_38_fu_3702_p2);

assign xor_ln45_94_fu_3152_p2 = (z1_29_fu_3064_p3 ^ z0_28_fu_2958_p3);

assign xor_ln45_95_fu_3158_p2 = (z2_182_fu_3130_p3 ^ tmp_13_fu_3144_p3);

assign xor_ln45_98_fu_3528_p2 = (z1_33_fu_3440_p3 ^ z0_33_fu_3334_p3);

assign xor_ln45_99_fu_3534_p2 = (z2_183_fu_3506_p3 ^ tmp_14_fu_3520_p3);

assign xor_ln45_9_fu_834_p2 = (z2_174_fu_794_p3 ^ z0_1_fu_622_p3);

assign xor_ln45_fu_610_p2 = (z1_fu_598_p2 ^ z0_fu_580_p2);

assign xor_ln59_13_fu_4590_p2 = (a1_sqr_30_fu_4512_p4 ^ a0_sqr_7_fu_4344_p4);

assign xor_ln59_14_fu_4596_p2 = (xor_ln59_9_fu_4406_p2 ^ tmp_23_fu_4492_p3);

assign xor_ln59_16_fu_6646_p2 = (a1_sqr_31_fu_6639_p3 ^ a0_sqr_16_fu_6628_p3);

assign xor_ln59_19_fu_6701_p2 = (a1_sqr_33_fu_6682_p3 ^ a0_sqr_18_fu_6652_p3);

assign xor_ln59_21_fu_7244_p2 = (a1_sqr_34_fu_7236_p3 ^ a0_sqr_23_fu_7228_p3);

assign xor_ln59_2_fu_4216_p2 = (a1_sqr_fu_4208_p3 ^ a0_sqr_1_fu_4178_p3);

assign xor_ln59_6_fu_4338_p2 = (a1_sqr_26_fu_4316_p3 ^ a0_sqr_3_fu_4232_p3);

assign xor_ln59_9_fu_4406_p2 = (a1_sqr_27_fu_4398_p3 ^ a0_sqr_9_fu_4368_p3);

assign xor_ln68_1_fu_4698_p2 = (tmp_104_fu_4582_p3 ^ tmp_103_fu_4574_p3);

assign xor_ln68_3_fu_4710_p2 = (xor_ln68_fu_4692_p2 ^ xor_ln68_1_fu_4698_p2);

assign xor_ln68_fu_4692_p2 = (tmp_99_fu_4038_p3 ^ tmp_102_fu_4068_p3);

assign xor_ln70_10_fu_4880_p2 = (xor_ln45_89_fu_3632_p2 ^ a0_69_fu_3804_p2);

assign xor_ln70_11_fu_4886_p2 = (xor_ln45_69_fu_2952_p2 ^ a0_57_fu_3124_p2);

assign xor_ln70_12_fu_4892_p2 = (xor_ln70_11_fu_4886_p2 ^ xor_ln70_10_fu_4880_p2);

assign xor_ln70_13_fu_4898_p2 = (xor_ln45_1_fu_616_p2 ^ a0_fu_788_p2);

assign xor_ln70_14_fu_4904_p2 = (xor_ln45_21_fu_1296_p2 ^ a0_23_fu_1468_p2);

assign xor_ln70_15_fu_4910_p2 = (xor_ln70_14_fu_4904_p2 ^ xor_ln70_13_fu_4898_p2);

assign xor_ln70_16_fu_4916_p2 = (xor_ln70_15_fu_4910_p2 ^ xor_ln70_12_fu_4892_p2);

assign xor_ln70_18_fu_4928_p2 = (xor_ln59_2_fu_4216_p2 ^ a0_86_fu_4300_p2);

assign xor_ln70_1_fu_446_p2 = (trunc_ln68_1_fu_172_p1 ^ tmp_98_fu_432_p3);

assign xor_ln70_20_fu_4934_p2 = (xor_ln70_18_fu_4928_p2 ^ xor_ln28_33_fu_4562_p2);

assign xor_ln70_21_fu_4940_p2 = (xor_ln45_41_fu_1610_p2 ^ xor_ln45_131_fu_3946_p2);

assign xor_ln70_23_fu_4952_p2 = (xor_ln59_6_fu_4338_p2 ^ a0_96_fu_4506_p2);

assign xor_ln70_24_fu_4958_p2 = (xor_ln45_33_fu_1598_p2 ^ a0_73_fu_3934_p2);

assign xor_ln70_27_fu_4984_p2 = (xor_ln68_3_fu_4710_p2 ^ tmp_111_fu_4970_p3);

assign xor_ln70_28_fu_6813_p2 = (b_198_fu_6624_p2 ^ a0_359_fu_6635_p2);

assign xor_ln70_29_fu_6819_p2 = (b_224_fu_6659_p2 ^ a0_361_reg_14151);

assign xor_ln70_2_fu_452_p2 = (trunc_ln68_2_fu_176_p1 ^ tmp_97_fu_424_p3);

assign xor_ln70_30_fu_6824_p2 = (xor_ln70_29_fu_6819_p2 ^ xor_ln70_28_fu_6813_p2);

assign xor_ln70_31_fu_6830_p2 = (xor_ln45_127_fu_6378_p2 ^ a0_128_fu_6474_p2);

assign xor_ln70_32_fu_6836_p2 = (xor_ln45_107_fu_5996_p2 ^ a0_111_fu_6092_p2);

assign xor_ln70_33_fu_6842_p2 = (xor_ln70_32_fu_6836_p2 ^ xor_ln70_31_fu_6830_p2);

assign xor_ln70_35_fu_6854_p2 = (xor_ln59_16_fu_6646_p2 ^ a0_138_fu_6676_p2);

assign xor_ln70_36_fu_6860_p2 = (xor_ln45_115_fu_6138_p2 ^ a0_129_fu_6520_p2);

assign xor_ln70_3_fu_458_p2 = (trunc_ln68_3_fu_180_p1 ^ tmp_96_fu_416_p3);

assign xor_ln70_4_fu_4844_p2 = (b_238_fu_4172_p2 ^ a0_331_fu_4202_p2);

assign xor_ln70_5_fu_4850_p2 = (xor_ln70_fu_4838_p2 ^ xor_ln70_4_fu_4844_p2);

assign xor_ln70_6_fu_4856_p2 = (b_344_fu_4446_p2 ^ a0_339_fu_260_p2);

assign xor_ln70_7_fu_4862_p2 = (b_318_fu_4362_p2 ^ a0_337_fu_4392_p2);

assign xor_ln70_8_fu_4868_p2 = (xor_ln70_7_fu_4862_p2 ^ xor_ln70_6_fu_4856_p2);

assign xor_ln70_9_fu_4874_p2 = (xor_ln70_8_fu_4868_p2 ^ xor_ln70_5_fu_4850_p2);

assign xor_ln70_fu_4838_p2 = (b_264_fu_4256_p2 ^ a0_334_fu_4286_p2);

assign xor_ln71_1_fu_4674_p2 = (tmp_110_fu_4656_p5 ^ tmp_109_fu_4648_p3);

assign xor_ln71_2_fu_4680_p2 = (tmp_108_fu_4640_p3 ^ tmp_107_fu_4632_p3);

assign xor_ln71_3_fu_4686_p2 = (tmp_106_fu_4622_p4 ^ tmp_105_fu_4614_p3);

assign xor_ln71_4_fu_6737_p2 = (tmp_113_fu_6724_p3 ^ tmp_112_fu_6716_p3);

assign xor_ln73_1_fu_9267_p2 = (xor_ln45_260_fu_8680_p2 ^ xor_ln45_259_fu_8674_p2);

assign xor_ln73_fu_9261_p2 = (xor_ln45_185_fu_8115_p2 ^ a0_201_fu_8608_p2);

assign z0_100_fu_9597_p3 = {{xor_ln45_254_fu_9585_p2}, {xor_ln45_255_fu_9591_p2}};

assign z0_101_fu_9638_p2 = (b0_71_fu_9633_p2 & a0_401_fu_9619_p2);

assign z0_102_fu_9694_p2 = (b0_72_reg_14460_pp0_iter1_reg & a0_402_fu_9605_p3);

assign z0_103_fu_9804_p2 = (a0_404_fu_9515_p1 & a0_332_reg_14062_pp0_iter1_reg);

assign z0_104_fu_9837_p3 = {{xor_ln45_264_fu_9825_p2}, {xor_ln45_265_fu_9831_p2}};

assign z0_105_fu_9877_p2 = (b0_74_fu_9873_p2 & a0_405_fu_9859_p2);

assign z0_106_fu_9933_p2 = (a0_406_fu_9845_p3 & a0_333_reg_14079_pp0_iter1_reg);

assign z0_107_fu_10084_p3 = {{xor_ln45_276_fu_10072_p2}, {xor_ln45_277_fu_10078_p2}};

assign z0_108_fu_10174_p2 = (b0_77_fu_10170_p2 & a0_409_fu_10156_p2);

assign z0_109_fu_10214_p3 = {{xor_ln45_278_fu_10202_p2}, {xor_ln45_279_fu_10208_p2}};

assign z0_10_fu_1302_p3 = {{xor_ln45_20_fu_1290_p2}, {xor_ln45_21_fu_1296_p2}};

assign z0_110_fu_10255_p2 = (b0_78_fu_10250_p2 & a0_410_fu_10236_p2);

assign z0_111_fu_10311_p2 = (b0_79_reg_14491_pp0_iter1_reg & a0_411_fu_10222_p3);

assign z0_112_fu_10395_p3 = {{xor_ln45_286_fu_10383_p2}, {xor_ln45_287_fu_10389_p2}};

assign z0_113_fu_10462_p2 = (b0_81_fu_10457_p2 & a0_413_fu_10443_p2);

assign z0_114_fu_10502_p3 = {{xor_ln45_288_fu_10490_p2}, {xor_ln45_289_fu_10496_p2}};

assign z0_115_fu_10543_p2 = (b0_82_fu_10538_p2 & a0_414_fu_10524_p2);

assign z0_116_fu_10599_p2 = (b0_83_reg_14524_pp0_iter1_reg & a0_415_fu_10510_p3);

assign z0_117_fu_10709_p2 = (b0_85_reg_14510_pp0_iter1_reg & a0_417_fu_10403_p3);

assign z0_118_fu_10747_p3 = {{xor_ln45_298_fu_10735_p2}, {xor_ln45_299_fu_10741_p2}};

assign z0_119_fu_10787_p2 = (b0_86_fu_10783_p2 & a0_418_fu_10769_p2);

assign z0_11_fu_1366_p2 = (b0_12_fu_1352_p2 & a0_301_fu_1338_p2);

assign z0_120_fu_10843_p2 = (b0_87_reg_14549_pp0_iter1_reg & a0_419_fu_10755_p3);

assign z0_121_fu_11025_p2 = (a0_422_fu_10092_p1 & a0_335_reg_13615_pp0_iter1_reg);

assign z0_122_fu_11058_p3 = {{xor_ln45_312_fu_11046_p2}, {xor_ln45_313_fu_11052_p2}};

assign z0_123_fu_11098_p2 = (b0_89_fu_11094_p2 & a0_423_fu_11080_p2);

assign z0_124_fu_11154_p2 = (a0_424_fu_11066_p3 & a0_336_reg_14105_pp0_iter1_reg);

assign z0_125_fu_11233_p3 = {{xor_ln45_320_fu_11221_p2}, {xor_ln45_321_fu_11227_p2}};

assign z0_126_fu_11285_p2 = (b0_91_fu_11281_p2 & a0_426_fu_11267_p2);

assign z0_127_fu_11325_p3 = {{xor_ln45_322_fu_11313_p2}, {xor_ln45_323_fu_11319_p2}};

assign z0_128_fu_11366_p2 = (b0_92_fu_11361_p2 & a0_427_fu_11347_p2);

assign z0_129_fu_11422_p2 = (b0_93_reg_14580_pp0_iter1_reg & a0_428_fu_11333_p3);

assign z0_12_fu_1432_p2 = (b0_13_fu_1324_p3 & a0_302_fu_1310_p3);

assign z0_130_fu_11532_p2 = (a0_430_fu_11241_p1 & a0_338_reg_14121_pp0_iter1_reg);

assign z0_131_fu_11565_p3 = {{xor_ln45_332_fu_11553_p2}, {xor_ln45_333_fu_11559_p2}};

assign z0_132_fu_11605_p2 = (b0_94_fu_11601_p2 & a0_431_fu_11587_p2);

assign z0_133_fu_11661_p2 = (a0_432_fu_11573_p3 & a0_288_reg_13599_pp0_iter1_reg);

assign z0_134_fu_11916_p2 = (b0_3_reg_13623_pp0_iter1_reg & a0_396_fu_9233_p2);

assign z0_135_fu_11943_p3 = {{xor_ln45_350_fu_11931_p2}, {xor_ln45_351_fu_11937_p2}};

assign z0_136_fu_11951_p2 = (b0_4_reg_13643_pp0_iter1_reg & a0_397_fu_9354_p2);

assign z0_137_fu_11986_p2 = (b0_5_reg_13638_pp0_iter1_reg & a0_398_fu_9340_p3);

assign z0_138_fu_12059_p3 = {{xor_ln45_358_fu_12047_p2}, {xor_ln45_359_fu_12053_p2}};

assign z0_139_fu_12067_p2 = (b0_7_reg_13673_pp0_iter1_reg & a0_400_fu_9539_p2);

assign z0_13_fu_1616_p3 = {{xor_ln45_32_fu_1592_p2}, {xor_ln45_33_fu_1598_p2}};

assign z0_140_fu_12094_p3 = {{xor_ln45_360_fu_12082_p2}, {xor_ln45_361_fu_12088_p2}};

assign z0_141_fu_12102_p2 = (b0_8_reg_13693_pp0_iter1_reg & a0_401_fu_9619_p2);

assign z0_142_fu_12137_p2 = (b0_9_reg_13688_pp0_iter1_reg & a0_402_fu_9605_p3);

assign z0_143_fu_12218_p2 = (b0_11_reg_13668_pp0_iter1_reg & a0_404_fu_9515_p1);

assign z0_144_fu_12245_p3 = {{xor_ln45_370_fu_12233_p2}, {xor_ln45_371_fu_12239_p2}};

assign z0_145_fu_12253_p2 = (b0_12_reg_13733_pp0_iter1_reg & a0_405_fu_9859_p2);

assign z0_146_fu_12288_p2 = (b0_13_reg_13728_pp0_iter1_reg & a0_406_fu_9845_p3);

assign z0_147_fu_12433_p3 = {{xor_ln45_382_fu_12421_p2}, {xor_ln45_383_fu_12427_p2}};

assign z0_148_fu_12441_p2 = (b0_16_reg_13763_pp0_iter1_reg & a0_409_fu_10156_p2);

assign z0_149_fu_12468_p3 = {{xor_ln45_384_fu_12456_p2}, {xor_ln45_385_fu_12462_p2}};

assign z0_14_fu_1816_p2 = (b0_16_fu_1802_p2 & a0_305_fu_1788_p2);

assign z0_150_fu_12476_p2 = (b0_17_reg_13783_pp0_iter1_reg & a0_410_fu_10236_p2);

assign z0_151_fu_12511_p2 = (b0_18_reg_13778_pp0_iter1_reg & a0_411_fu_10222_p3);

assign z0_152_fu_12584_p3 = {{xor_ln45_392_fu_12572_p2}, {xor_ln45_393_fu_12578_p2}};

assign z0_153_fu_12592_p2 = (b0_20_reg_13813_pp0_iter1_reg & a0_413_fu_10443_p2);

assign z0_154_fu_12619_p3 = {{xor_ln45_394_fu_12607_p2}, {xor_ln45_395_fu_12613_p2}};

assign z0_155_fu_12627_p2 = (b0_21_reg_13833_pp0_iter1_reg & a0_414_fu_10524_p2);

assign z0_156_fu_12662_p2 = (b0_22_reg_13828_pp0_iter1_reg & a0_415_fu_10510_p3);

assign z0_157_fu_12743_p2 = (b0_24_reg_13808_pp0_iter1_reg & a0_417_fu_10403_p3);

assign z0_158_fu_12770_p3 = {{xor_ln45_404_fu_12758_p2}, {xor_ln45_405_fu_12764_p2}};

assign z0_159_fu_12778_p2 = (b0_25_reg_13873_pp0_iter1_reg & a0_418_fu_10769_p2);

assign z0_15_fu_1858_p3 = {{xor_ln45_34_fu_1846_p2}, {xor_ln45_35_fu_1852_p2}};

assign z0_160_fu_12813_p2 = (b0_26_reg_13868_pp0_iter1_reg & a0_419_fu_10755_p3);

assign z0_161_fu_12966_p2 = (b0_29_reg_13758_pp0_iter1_reg & a0_422_fu_10092_p1);

assign z0_162_fu_12993_p3 = {{xor_ln45_418_fu_12981_p2}, {xor_ln45_419_fu_12987_p2}};

assign z0_163_fu_13001_p2 = (b0_30_reg_13913_pp0_iter1_reg & a0_423_fu_11080_p2);

assign z0_164_fu_13036_p2 = (b0_31_reg_13908_pp0_iter1_reg & a0_424_fu_11066_p3);

assign z0_165_fu_13109_p3 = {{xor_ln45_426_fu_13097_p2}, {xor_ln45_427_fu_13103_p2}};

assign z0_166_fu_13117_p2 = (b0_33_reg_13943_pp0_iter1_reg & a0_426_fu_11267_p2);

assign z0_167_fu_13144_p3 = {{xor_ln45_428_fu_13132_p2}, {xor_ln45_429_fu_13138_p2}};

assign z0_168_fu_13152_p2 = (b0_34_reg_13963_pp0_iter1_reg & a0_427_fu_11347_p2);

assign z0_169_fu_13187_p2 = (b0_35_reg_13958_pp0_iter1_reg & a0_428_fu_11333_p3);

assign z0_16_fu_1922_p2 = (b0_17_fu_1908_p2 & a0_306_fu_1894_p2);

assign z0_170_fu_13268_p2 = (b0_37_reg_13938_pp0_iter1_reg & a0_430_fu_11241_p1);

assign z0_171_fu_13295_p3 = {{xor_ln45_438_fu_13283_p2}, {xor_ln45_439_fu_13289_p2}};

assign z0_172_fu_13303_p2 = (b0_38_reg_14003_pp0_iter1_reg & a0_431_fu_11587_p2);

assign z0_173_fu_13338_p2 = (b0_39_reg_13998_pp0_iter1_reg & a0_432_fu_11573_p3);

assign z0_17_fu_1988_p2 = (b0_18_fu_1880_p3 & a0_307_fu_1866_p3);

assign z0_18_fu_2076_p3 = {{xor_ln45_42_fu_2064_p2}, {xor_ln45_43_fu_2070_p2}};

assign z0_19_fu_2192_p2 = (b0_20_fu_2178_p2 & a0_309_fu_2164_p2);

assign z0_1_fu_622_p3 = {{xor_ln45_fu_610_p2}, {xor_ln45_1_fu_616_p2}};

assign z0_20_fu_2234_p3 = {{xor_ln45_44_fu_2222_p2}, {xor_ln45_45_fu_2228_p2}};

assign z0_21_fu_2298_p2 = (b0_21_fu_2284_p2 & a0_310_fu_2270_p2);

assign z0_22_fu_2364_p2 = (b0_22_fu_2256_p3 & a0_311_fu_2242_p3);

assign z0_23_fu_2496_p2 = (b0_24_fu_2108_p3 & a0_313_fu_2084_p3);

assign z0_24_fu_2538_p3 = {{xor_ln45_54_fu_2526_p2}, {xor_ln45_55_fu_2532_p2}};

assign z0_25_fu_2602_p2 = (b0_25_fu_2588_p2 & a0_314_fu_2574_p2);

assign z0_26_fu_2668_p2 = (b0_26_fu_2560_p3 & a0_315_fu_2546_p3);

assign z0_27_fu_2916_p2 = (b0_29_fu_1674_p3 & a0_318_fu_1624_p3);

assign z0_28_fu_2958_p3 = {{xor_ln45_68_fu_2946_p2}, {xor_ln45_69_fu_2952_p2}};

assign z0_29_fu_3022_p2 = (b0_30_fu_3008_p2 & a0_319_fu_2994_p2);

assign z0_2_fu_686_p2 = (b0_4_fu_672_p2 & a0_293_fu_658_p2);

assign z0_30_fu_3088_p2 = (b0_31_fu_2980_p3 & a0_320_fu_2966_p3);

assign z0_31_fu_3176_p3 = {{xor_ln45_76_fu_3164_p2}, {xor_ln45_77_fu_3170_p2}};

assign z0_32_fu_3292_p2 = (b0_33_fu_3278_p2 & a0_322_fu_3264_p2);

assign z0_33_fu_3334_p3 = {{xor_ln45_78_fu_3322_p2}, {xor_ln45_79_fu_3328_p2}};

assign z0_34_fu_3398_p2 = (b0_34_fu_3384_p2 & a0_323_fu_3370_p2);

assign z0_35_fu_3464_p2 = (b0_35_fu_3356_p3 & a0_324_fu_3342_p3);

assign z0_36_fu_3596_p2 = (b0_37_fu_3208_p3 & a0_326_fu_3184_p3);

assign z0_37_fu_3638_p3 = {{xor_ln45_88_fu_3626_p2}, {xor_ln45_89_fu_3632_p2}};

assign z0_38_fu_3702_p2 = (b0_38_fu_3688_p2 & a0_327_fu_3674_p2);

assign z0_39_fu_3768_p2 = (b0_39_fu_3660_p3 & a0_328_fu_3646_p3);

assign z0_3_fu_752_p2 = (b0_5_fu_644_p3 & a0_294_fu_630_p3);

assign z0_40_fu_5968_p2 = (b0_42_reg_14181 & a0_346_reg_14167);

assign z0_41_fu_6002_p3 = {{xor_ln45_106_fu_5990_p2}, {xor_ln45_107_fu_5996_p2}};

assign z0_42_fu_6018_p2 = (b0_43_fu_6014_p2 & a0_347_fu_6010_p2);

assign z0_43_fu_6064_p2 = (b0_44_reg_14204 & a0_348_reg_14197);

assign z0_44_fu_6144_p3 = {{xor_ln45_114_fu_6132_p2}, {xor_ln45_115_fu_6138_p2}};

assign z0_45_fu_6160_p2 = (b0_46_fu_6156_p2 & a0_350_fu_6152_p2);

assign z0_46_fu_6198_p3 = {{xor_ln45_116_fu_6186_p2}, {xor_ln45_117_fu_6192_p2}};

assign z0_47_fu_6216_p2 = (b0_47_fu_6211_p2 & a0_351_fu_6206_p2);

assign z0_48_fu_6262_p2 = (b0_48_reg_14275 & a0_352_reg_14268);

assign z0_49_fu_6350_p2 = (b0_50_reg_14246 & a0_354_reg_14238);

assign z0_4_fu_840_p3 = {{xor_ln45_8_fu_828_p2}, {xor_ln45_9_fu_834_p2}};

assign z0_50_fu_6384_p3 = {{xor_ln45_126_fu_6372_p2}, {xor_ln45_127_fu_6378_p2}};

assign z0_51_fu_6400_p2 = (b0_51_fu_6396_p2 & a0_355_fu_6392_p2);

assign z0_52_fu_6446_p2 = (b0_52_reg_14329 & a0_356_reg_14322);

assign z0_53_fu_6926_p2 = (b0_54_fu_6912_p2 & a0_366_fu_6848_p2);

assign z0_54_fu_6968_p3 = {{xor_ln45_140_fu_6956_p2}, {xor_ln45_141_fu_6962_p2}};

assign z0_55_fu_7032_p2 = (b0_55_fu_7018_p2 & a0_367_fu_7004_p2);

assign z0_56_fu_7098_p2 = (b0_56_fu_6990_p3 & a0_368_fu_6976_p3);

assign z0_57_fu_7378_p2 = (b0_57_fu_7356_p2 & a0_373_fu_7308_p2);

assign z0_58_fu_7486_p2 = (a0_375_fu_7480_p2 & a0_372_fu_7320_p3);

assign z0_59_fu_7522_p2 = (b0_57_fu_7356_p2 & a0_375_fu_7480_p2);

assign z0_5_fu_956_p2 = (b0_7_fu_942_p2 & a0_296_fu_928_p2);

assign z0_60_fu_7590_p2 = (a0_377_reg_14784 & a0_369_reg_14746);

assign z0_61_fu_7614_p3 = {{xor_ln45_156_fu_7602_p2}, {xor_ln45_157_fu_7608_p2}};

assign z0_62_fu_7644_p2 = (b0_58_fu_7640_p2 & a0_378_fu_7628_p2);

assign z0_63_fu_7692_p2 = (a0_379_reg_14769 & a0_364_reg_14685);

assign z0_64_fu_7762_p2 = (b0_54_reg_14701 & a0_377_reg_14784);

assign z0_65_fu_7786_p3 = {{xor_ln45_166_fu_7774_p2}, {xor_ln45_167_fu_7780_p2}};

assign z0_66_fu_7794_p2 = (b0_55_reg_14721 & a0_378_fu_7628_p2);

assign z0_67_fu_7829_p2 = (b0_56_reg_14716 & a0_379_reg_14769);

assign z0_68_fu_7923_p2 = (a0_382_fu_7893_p2 & a0_357_reg_14363_pp0_iter1_reg);

assign z0_69_fu_7956_p3 = {{xor_ln45_176_fu_7944_p2}, {xor_ln45_177_fu_7950_p2}};

assign z0_6_fu_998_p3 = {{xor_ln45_10_fu_986_p2}, {xor_ln45_11_fu_992_p2}};

assign z0_70_fu_7986_p2 = (b0_60_fu_7982_p2 & a0_383_fu_7968_p2);

assign z0_71_fu_8042_p2 = (a0_384_fu_7964_p1 & a0_358_reg_14378_pp0_iter1_reg);

assign z0_72_fu_8121_p3 = {{xor_ln45_184_fu_8109_p2}, {xor_ln45_185_fu_8115_p2}};

assign z0_73_fu_8173_p2 = (b0_62_fu_8169_p2 & a0_386_fu_8155_p2);

assign z0_74_fu_8213_p3 = {{xor_ln45_186_fu_8201_p2}, {xor_ln45_187_fu_8207_p2}};

assign z0_75_fu_8254_p2 = (b0_63_fu_8249_p2 & a0_387_fu_8235_p2);

assign z0_76_fu_8310_p2 = (b0_64_reg_14423_pp0_iter1_reg & a0_388_fu_8221_p3);

assign z0_77_fu_8410_p2 = (a0_390_fu_8129_p1 & a0_360_reg_14159_pp0_iter1_reg);

assign z0_78_fu_8443_p3 = {{xor_ln45_196_fu_8431_p2}, {xor_ln45_197_fu_8437_p2}};

assign z0_79_fu_8479_p2 = (b0_65_fu_8475_p2 & a0_391_fu_8461_p2);

assign z0_7_fu_1062_p2 = (b0_8_fu_1048_p2 & a0_297_fu_1034_p2);

assign z0_80_fu_8535_p2 = (a0_392_fu_8451_p1 & a0_343_reg_14138_pp0_iter1_reg);

assign z0_81_fu_8698_p2 = (b0_42_reg_14181_pp0_iter1_reg & a0_382_fu_7893_p2);

assign z0_82_fu_8725_p3 = {{xor_ln45_210_fu_8713_p2}, {xor_ln45_211_fu_8719_p2}};

assign z0_83_fu_8733_p2 = (b0_43_reg_14610 & a0_383_fu_7968_p2);

assign z0_84_fu_8768_p2 = (b0_44_reg_14204_pp0_iter1_reg & a0_384_fu_7964_p1);

assign z0_85_fu_8841_p3 = {{xor_ln45_218_fu_8829_p2}, {xor_ln45_219_fu_8835_p2}};

assign z0_86_fu_8849_p2 = (b0_46_reg_14625 & a0_386_fu_8155_p2);

assign z0_87_fu_8876_p3 = {{xor_ln45_220_fu_8864_p2}, {xor_ln45_221_fu_8870_p2}};

assign z0_88_fu_8884_p2 = (b0_47_reg_14635 & a0_387_fu_8235_p2);

assign z0_89_fu_8919_p2 = (b0_48_reg_14275_pp0_iter1_reg & a0_388_fu_8221_p3);

assign z0_8_fu_1128_p2 = (b0_9_fu_1020_p3 & a0_298_fu_1006_p3);

assign z0_90_fu_9000_p2 = (b0_50_reg_14246_pp0_iter1_reg & a0_390_fu_8129_p1);

assign z0_91_fu_9027_p3 = {{xor_ln45_230_fu_9015_p2}, {xor_ln45_231_fu_9021_p2}};

assign z0_92_fu_9035_p2 = (b0_51_reg_14655 & a0_391_fu_8461_p2);

assign z0_93_fu_9070_p2 = (b0_52_reg_14329_pp0_iter1_reg & a0_392_fu_8451_p1);

assign z0_94_fu_9299_p2 = (a0_396_fu_9233_p2 & a0_329_reg_14028_pp0_iter1_reg);

assign z0_95_fu_9332_p3 = {{xor_ln45_244_fu_9320_p2}, {xor_ln45_245_fu_9326_p2}};

assign z0_96_fu_9372_p2 = (b0_68_fu_9368_p2 & a0_397_fu_9354_p2);

assign z0_97_fu_9428_p2 = (a0_398_fu_9340_p3 & a0_330_reg_14046_pp0_iter1_reg);

assign z0_98_fu_9507_p3 = {{xor_ln45_252_fu_9495_p2}, {xor_ln45_253_fu_9501_p2}};

assign z0_99_fu_9557_p2 = (b0_70_fu_9553_p2 & a0_400_fu_9539_p2);

assign z0_9_fu_1260_p2 = (b0_11_fu_872_p3 & a0_300_fu_848_p3);

assign z0_fu_580_p2 = (b0_3_fu_566_p2 & a0_292_fu_396_p1);

assign z1_100_fu_9678_p3 = {{xor_ln45_256_fu_9666_p2}, {xor_ln45_257_fu_9672_p2}};

assign z1_101_fu_9709_p2 = (b_259_fu_9705_p2 & a_320_fu_9699_p2);

assign z1_102_fu_9778_p3 = {{xor_ln45_262_fu_9766_p2}, {xor_ln45_263_fu_9772_p2}};

assign z1_103_fu_9815_p2 = (b_264_reg_14074_pp0_iter1_reg & a_326_fu_9809_p2);

assign z1_104_fu_9894_p2 = (b_268_fu_9889_p2 & a_330_fu_9883_p2);

assign z1_105_fu_9917_p3 = {{xor_ln45_266_fu_9905_p2}, {xor_ln45_267_fu_9911_p2}};

assign z1_106_fu_9944_p2 = (a_334_fu_9938_p2 & a0_334_reg_14090_pp0_iter1_reg);

assign z1_107_fu_10191_p2 = (b_278_fu_10186_p2 & a_343_fu_10180_p2);

assign z1_108_fu_10272_p2 = (b_282_fu_10267_p2 & a_347_fu_10261_p2);

assign z1_109_fu_10295_p3 = {{xor_ln45_280_fu_10283_p2}, {xor_ln45_281_fu_10289_p2}};

assign z1_10_fu_1384_p2 = (b_35_fu_1378_p2 & a_41_fu_1372_p2);

assign z1_110_fu_10326_p2 = (b_286_fu_10322_p2 & a_351_fu_10316_p2);

assign z1_111_fu_10479_p2 = (b_291_fu_10474_p2 & a_357_fu_10468_p2);

assign z1_112_fu_10560_p2 = (b_295_fu_10555_p2 & a_361_fu_10549_p2);

assign z1_113_fu_10583_p3 = {{xor_ln45_290_fu_10571_p2}, {xor_ln45_291_fu_10577_p2}};

assign z1_114_fu_10614_p2 = (b_299_fu_10610_p2 & a_365_fu_10604_p2);

assign z1_115_fu_10683_p3 = {{xor_ln45_296_fu_10671_p2}, {xor_ln45_297_fu_10677_p2}};

assign z1_116_fu_10724_p2 = (b_304_fu_10720_p2 & a_371_fu_10714_p2);

assign z1_117_fu_10804_p2 = (b_308_fu_10799_p2 & a_375_fu_10793_p2);

assign z1_118_fu_10827_p3 = {{xor_ln45_300_fu_10815_p2}, {xor_ln45_301_fu_10821_p2}};

assign z1_119_fu_10858_p2 = (b_312_fu_10854_p2 & a_379_fu_10848_p2);

assign z1_11_fu_1408_p3 = {{xor_ln45_22_fu_1396_p2}, {xor_ln45_23_fu_1402_p2}};

assign z1_120_fu_10999_p3 = {{xor_ln45_310_fu_10987_p2}, {xor_ln45_311_fu_10993_p2}};

assign z1_121_fu_11036_p2 = (b_318_reg_14100_pp0_iter1_reg & a_388_fu_11030_p2);

assign z1_122_fu_11115_p2 = (b_322_fu_11110_p2 & a_392_fu_11104_p2);

assign z1_123_fu_11138_p3 = {{xor_ln45_314_fu_11126_p2}, {xor_ln45_315_fu_11132_p2}};

assign z1_124_fu_11165_p2 = (a_396_fu_11159_p2 & a0_337_reg_14116_pp0_iter1_reg);

assign z1_125_fu_11302_p2 = (b_331_fu_11297_p2 & a_402_fu_11291_p2);

assign z1_126_fu_11383_p2 = (b_335_fu_11378_p2 & a_406_fu_11372_p2);

assign z1_127_fu_11406_p3 = {{xor_ln45_324_fu_11394_p2}, {xor_ln45_325_fu_11400_p2}};

assign z1_128_fu_11437_p2 = (b_339_fu_11433_p2 & a_410_fu_11427_p2);

assign z1_129_fu_11506_p3 = {{xor_ln45_330_fu_11494_p2}, {xor_ln45_331_fu_11500_p2}};

assign z1_12_fu_1450_p2 = (b_39_fu_1444_p2 & a_45_fu_1438_p2);

assign z1_130_fu_11543_p2 = (b_344_reg_14133_pp0_iter1_reg & a_416_fu_11537_p2);

assign z1_131_fu_11622_p2 = (b_348_fu_11617_p2 & a_420_fu_11611_p2);

assign z1_132_fu_11645_p3 = {{xor_ln45_334_fu_11633_p2}, {xor_ln45_335_fu_11639_p2}};

assign z1_133_fu_11672_p2 = (a_424_fu_11666_p2 & a0_339_reg_13610_pp0_iter1_reg);

assign z1_134_fu_11921_p2 = (b_5_reg_13633_pp0_iter1_reg & a_298_fu_9304_p2);

assign z1_135_fu_11956_p2 = (b_9_reg_13653_pp0_iter1_reg & a_302_fu_9378_p2);

assign z1_136_fu_11978_p3 = {{xor_ln45_352_fu_11966_p2}, {xor_ln45_353_fu_11972_p2}};

assign z1_137_fu_11991_p2 = (b_13_reg_13663_pp0_iter1_reg & a_306_fu_9433_p2);

assign z1_138_fu_12072_p2 = (b_18_reg_13683_pp0_iter1_reg & a_312_fu_9563_p2);

assign z1_139_fu_12107_p2 = (b_22_reg_13703_pp0_iter1_reg & a_316_fu_9644_p2);

assign z1_13_fu_1834_p2 = (b_45_fu_1828_p2 & a_54_fu_1822_p2);

assign z1_140_fu_12129_p3 = {{xor_ln45_362_fu_12117_p2}, {xor_ln45_363_fu_12123_p2}};

assign z1_141_fu_12142_p2 = (b_26_reg_13713_pp0_iter1_reg & a_320_fu_9699_p2);

assign z1_142_fu_12210_p3 = {{xor_ln45_368_fu_12198_p2}, {xor_ln45_369_fu_12204_p2}};

assign z1_143_fu_12223_p2 = (b_31_reg_13723_pp0_iter1_reg & a_326_fu_9809_p2);

assign z1_144_fu_12258_p2 = (b_35_reg_13743_pp0_iter1_reg & a_330_fu_9883_p2);

assign z1_145_fu_12280_p3 = {{xor_ln45_372_fu_12268_p2}, {xor_ln45_373_fu_12274_p2}};

assign z1_146_fu_12293_p2 = (b_39_reg_13753_pp0_iter1_reg & a_334_fu_9938_p2);

assign z1_147_fu_12446_p2 = (b_45_reg_13773_pp0_iter1_reg & a_343_fu_10180_p2);

assign z1_148_fu_12481_p2 = (b_49_reg_13793_pp0_iter1_reg & a_347_fu_10261_p2);

assign z1_149_fu_12503_p3 = {{xor_ln45_386_fu_12491_p2}, {xor_ln45_387_fu_12497_p2}};

assign z1_14_fu_1940_p2 = (b_49_fu_1934_p2 & a_58_fu_1928_p2);

assign z1_150_fu_12516_p2 = (b_53_reg_13803_pp0_iter1_reg & a_351_fu_10316_p2);

assign z1_151_fu_12597_p2 = (b_58_reg_13823_pp0_iter1_reg & a_357_fu_10468_p2);

assign z1_152_fu_12632_p2 = (b_62_reg_13843_pp0_iter1_reg & a_361_fu_10549_p2);

assign z1_153_fu_12654_p3 = {{xor_ln45_396_fu_12642_p2}, {xor_ln45_397_fu_12648_p2}};

assign z1_154_fu_12667_p2 = (b_66_reg_13853_pp0_iter1_reg & a_365_fu_10604_p2);

assign z1_155_fu_12735_p3 = {{xor_ln45_402_fu_12723_p2}, {xor_ln45_403_fu_12729_p2}};

assign z1_156_fu_12748_p2 = (b_71_reg_13863_pp0_iter1_reg & a_371_fu_10714_p2);

assign z1_157_fu_12783_p2 = (b_75_reg_13883_pp0_iter1_reg & a_375_fu_10793_p2);

assign z1_158_fu_12805_p3 = {{xor_ln45_406_fu_12793_p2}, {xor_ln45_407_fu_12799_p2}};

assign z1_159_fu_12818_p2 = (b_79_reg_13893_pp0_iter1_reg & a_379_fu_10848_p2);

assign z1_15_fu_1964_p3 = {{xor_ln45_36_fu_1952_p2}, {xor_ln45_37_fu_1958_p2}};

assign z1_160_fu_12958_p3 = {{xor_ln45_416_fu_12946_p2}, {xor_ln45_417_fu_12952_p2}};

assign z1_161_fu_12971_p2 = (b_85_reg_13903_pp0_iter1_reg & a_388_fu_11030_p2);

assign z1_162_fu_13006_p2 = (b_89_reg_13923_pp0_iter1_reg & a_392_fu_11104_p2);

assign z1_163_fu_13028_p3 = {{xor_ln45_420_fu_13016_p2}, {xor_ln45_421_fu_13022_p2}};

assign z1_164_fu_13041_p2 = (b_93_reg_13933_pp0_iter1_reg & a_396_fu_11159_p2);

assign z1_165_fu_13122_p2 = (b_98_reg_13953_pp0_iter1_reg & a_402_fu_11291_p2);

assign z1_166_fu_13157_p2 = (b_102_reg_13973_pp0_iter1_reg & a_406_fu_11372_p2);

assign z1_167_fu_13179_p3 = {{xor_ln45_430_fu_13167_p2}, {xor_ln45_431_fu_13173_p2}};

assign z1_168_fu_13192_p2 = (b_106_reg_13983_pp0_iter1_reg & a_410_fu_11427_p2);

assign z1_169_fu_13260_p3 = {{xor_ln45_436_fu_13248_p2}, {xor_ln45_437_fu_13254_p2}};

assign z1_16_fu_2006_p2 = (b_53_fu_2000_p2 & a_62_fu_1994_p2);

assign z1_170_fu_13273_p2 = (b_111_reg_13993_pp0_iter1_reg & a_416_fu_11537_p2);

assign z1_171_fu_13308_p2 = (b_115_reg_14013_pp0_iter1_reg & a_420_fu_11611_p2);

assign z1_172_fu_13330_p3 = {{xor_ln45_440_fu_13318_p2}, {xor_ln45_441_fu_13324_p2}};

assign z1_173_fu_13343_p2 = (b_119_reg_14023_pp0_iter1_reg & a_424_fu_11666_p2);

assign z1_17_fu_2210_p2 = (b_58_fu_2204_p2 & a_68_fu_2198_p2);

assign z1_18_fu_2316_p2 = (b_62_fu_2310_p2 & a_72_fu_2304_p2);

assign z1_19_fu_2340_p3 = {{xor_ln45_46_fu_2328_p2}, {xor_ln45_47_fu_2334_p2}};

assign z1_1_fu_704_p2 = (b_9_fu_698_p2 & a_13_fu_692_p2);

assign z1_20_fu_2382_p2 = (b_66_fu_2376_p2 & a_76_fu_2370_p2);

assign z1_21_fu_2452_p3 = {{xor_ln45_52_fu_2440_p2}, {xor_ln45_53_fu_2446_p2}};

assign z1_22_fu_2514_p2 = (b_71_fu_2508_p2 & a_82_fu_2502_p2);

assign z1_23_fu_2620_p2 = (b_75_fu_2614_p2 & a_86_fu_2608_p2);

assign z1_24_fu_2644_p3 = {{xor_ln45_56_fu_2632_p2}, {xor_ln45_57_fu_2638_p2}};

assign z1_25_fu_2686_p2 = (b_79_fu_2680_p2 & a_90_fu_2674_p2);

assign z1_26_fu_2852_p3 = {{xor_ln45_66_fu_2828_p2}, {xor_ln45_67_fu_2834_p2}};

assign z1_27_fu_2934_p2 = (b_85_fu_2928_p2 & a_99_fu_2922_p2);

assign z1_28_fu_3040_p2 = (b_89_fu_3034_p2 & a_103_fu_3028_p2);

assign z1_29_fu_3064_p3 = {{xor_ln45_70_fu_3052_p2}, {xor_ln45_71_fu_3058_p2}};

assign z1_2_fu_728_p3 = {{xor_ln45_2_fu_716_p2}, {xor_ln45_3_fu_722_p2}};

assign z1_30_fu_3106_p2 = (b_93_fu_3100_p2 & a_107_fu_3094_p2);

assign z1_31_fu_3310_p2 = (b_98_fu_3304_p2 & a_113_fu_3298_p2);

assign z1_32_fu_3416_p2 = (b_102_fu_3410_p2 & a_117_fu_3404_p2);

assign z1_33_fu_3440_p3 = {{xor_ln45_80_fu_3428_p2}, {xor_ln45_81_fu_3434_p2}};

assign z1_34_fu_3482_p2 = (b_106_fu_3476_p2 & a_121_fu_3470_p2);

assign z1_35_fu_3552_p3 = {{xor_ln45_86_fu_3540_p2}, {xor_ln45_87_fu_3546_p2}};

assign z1_36_fu_3614_p2 = (b_111_fu_3608_p2 & a_127_fu_3602_p2);

assign z1_37_fu_3720_p2 = (b_115_fu_3714_p2 & a_131_fu_3708_p2);

assign z1_38_fu_3744_p3 = {{xor_ln45_90_fu_3732_p2}, {xor_ln45_91_fu_3738_p2}};

assign z1_39_fu_3786_p2 = (b_119_fu_3780_p2 & a_135_fu_3774_p2);

assign z1_3_fu_770_p2 = (b_13_fu_764_p2 & a_17_fu_758_p2);

assign z1_40_fu_5980_p2 = (b_125_fu_5976_p2 & a_159_fu_5972_p2);

assign z1_41_fu_6034_p2 = (b_129_fu_6029_p2 & a_163_fu_6024_p2);

assign z1_42_fu_6056_p3 = {{xor_ln45_108_fu_6044_p2}, {xor_ln45_109_fu_6050_p2}};

assign z1_43_fu_6076_p2 = (b_133_fu_6072_p2 & a_167_fu_6068_p2);

assign z1_44_fu_6176_p2 = (b_138_fu_6171_p2 & a_173_fu_6166_p2);

assign z1_45_fu_6232_p2 = (b_142_fu_6227_p2 & a_177_fu_6222_p2);

assign z1_46_fu_6254_p3 = {{xor_ln45_118_fu_6242_p2}, {xor_ln45_119_fu_6248_p2}};

assign z1_47_fu_6274_p2 = (b_146_fu_6270_p2 & a_181_fu_6266_p2);

assign z1_48_fu_6342_p3 = {{xor_ln45_124_fu_6330_p2}, {xor_ln45_125_fu_6336_p2}};

assign z1_49_fu_6362_p2 = (b_151_fu_6358_p2 & a_187_fu_6354_p2);

assign z1_4_fu_974_p2 = (b_18_fu_968_p2 & a_23_fu_962_p2);

assign z1_50_fu_6416_p2 = (b_155_fu_6411_p2 & a_191_fu_6406_p2);

assign z1_51_fu_6438_p3 = {{xor_ln45_128_fu_6426_p2}, {xor_ln45_129_fu_6432_p2}};

assign z1_52_fu_6458_p2 = (b_159_fu_6454_p2 & a_195_fu_6450_p2);

assign z1_53_fu_6944_p2 = (b_164_fu_6938_p2 & a_208_fu_6932_p2);

assign z1_54_fu_7050_p2 = (b_168_fu_7044_p2 & a_212_fu_7038_p2);

assign z1_55_fu_7074_p3 = {{xor_ln45_142_fu_7062_p2}, {xor_ln45_143_fu_7068_p2}};

assign z1_56_fu_7116_p2 = (b_172_fu_7110_p2 & a_216_fu_7104_p2);

assign z1_57_fu_7396_p2 = (b_176_fu_7390_p2 & a_223_fu_7384_p2);

assign z1_58_fu_7498_p2 = (b_181_fu_7336_p2 & a_229_fu_7492_p2);

assign z1_59_fu_7528_p2 = (b_176_fu_7390_p2 & a_229_fu_7492_p2);

assign z1_5_fu_1080_p2 = (b_22_fu_1074_p2 & a_27_fu_1068_p2);

assign z1_60_fu_7594_p2 = (b_185_reg_14757 & a_233_reg_14792);

assign z1_61_fu_7661_p2 = (b_189_fu_7656_p2 & a_237_fu_7650_p2);

assign z1_62_fu_7684_p3 = {{xor_ln45_158_fu_7672_p2}, {xor_ln45_159_fu_7678_p2}};

assign z1_63_fu_7696_p2 = (a_241_reg_14804 & a0_370_reg_14696);

assign z1_64_fu_7766_p2 = (b_164_reg_14711 & a_233_reg_14792);

assign z1_65_fu_7799_p2 = (b_168_reg_14731 & a_237_fu_7650_p2);

assign z1_66_fu_7821_p3 = {{xor_ln45_168_fu_7809_p2}, {xor_ln45_169_fu_7815_p2}};

assign z1_67_fu_7833_p2 = (b_172_reg_14741 & a_241_reg_14804);

assign z1_68_fu_7934_p2 = (b_198_reg_14670 & a_248_fu_7928_p2);

assign z1_69_fu_8003_p2 = (b_202_fu_7998_p2 & a_252_fu_7992_p2);

assign z1_6_fu_1104_p3 = {{xor_ln45_12_fu_1092_p2}, {xor_ln45_13_fu_1098_p2}};

assign z1_70_fu_8026_p3 = {{xor_ln45_178_fu_8014_p2}, {xor_ln45_179_fu_8020_p2}};

assign z1_71_fu_8053_p2 = (a_256_fu_8047_p2 & a0_359_reg_14675);

assign z1_72_fu_8190_p2 = (b_211_fu_8185_p2 & a_262_fu_8179_p2);

assign z1_73_fu_8271_p2 = (b_215_fu_8266_p2 & a_266_fu_8260_p2);

assign z1_74_fu_8294_p3 = {{xor_ln45_188_fu_8282_p2}, {xor_ln45_189_fu_8288_p2}};

assign z1_75_fu_8325_p2 = (b_219_fu_8321_p2 & a_270_fu_8315_p2);

assign z1_76_fu_8394_p3 = {{xor_ln45_194_fu_8382_p2}, {xor_ln45_195_fu_8388_p2}};

assign z1_77_fu_8421_p2 = (b_224_reg_14680 & a_276_fu_8415_p2);

assign z1_78_fu_8496_p2 = (b_228_fu_8491_p2 & a_280_fu_8485_p2);

assign z1_79_fu_8519_p3 = {{xor_ln45_198_fu_8507_p2}, {xor_ln45_199_fu_8513_p2}};

assign z1_7_fu_1146_p2 = (b_26_fu_1140_p2 & a_31_fu_1134_p2);

assign z1_80_fu_8546_p2 = (a_284_fu_8540_p2 & a0_361_reg_14151_pp0_iter1_reg);

assign z1_81_fu_8703_p2 = (b_125_reg_14605 & a_248_fu_7928_p2);

assign z1_82_fu_8738_p2 = (b_129_reg_14615 & a_252_fu_7992_p2);

assign z1_83_fu_8760_p3 = {{xor_ln45_212_fu_8748_p2}, {xor_ln45_213_fu_8754_p2}};

assign z1_84_fu_8773_p2 = (b_133_reg_14620 & a_256_fu_8047_p2);

assign z1_85_fu_8854_p2 = (b_138_reg_14630 & a_262_fu_8179_p2);

assign z1_86_fu_8889_p2 = (b_142_reg_14640 & a_266_fu_8260_p2);

assign z1_87_fu_8911_p3 = {{xor_ln45_222_fu_8899_p2}, {xor_ln45_223_fu_8905_p2}};

assign z1_88_fu_8924_p2 = (b_146_reg_14645 & a_270_fu_8315_p2);

assign z1_89_fu_8992_p3 = {{xor_ln45_228_fu_8980_p2}, {xor_ln45_229_fu_8986_p2}};

assign z1_8_fu_1216_p3 = {{xor_ln45_18_fu_1204_p2}, {xor_ln45_19_fu_1210_p2}};

assign z1_90_fu_9005_p2 = (b_151_reg_14650 & a_276_fu_8415_p2);

assign z1_91_fu_9040_p2 = (b_155_reg_14660 & a_280_fu_8485_p2);

assign z1_92_fu_9062_p3 = {{xor_ln45_232_fu_9050_p2}, {xor_ln45_233_fu_9056_p2}};

assign z1_93_fu_9075_p2 = (b_159_reg_14665 & a_284_fu_8540_p2);

assign z1_94_fu_9310_p2 = (b_238_reg_14041_pp0_iter1_reg & a_298_fu_9304_p2);

assign z1_95_fu_9389_p2 = (b_242_fu_9384_p2 & a_302_fu_9378_p2);

assign z1_96_fu_9412_p3 = {{xor_ln45_246_fu_9400_p2}, {xor_ln45_247_fu_9406_p2}};

assign z1_97_fu_9439_p2 = (a_306_fu_9433_p2 & a0_331_reg_14057_pp0_iter1_reg);

assign z1_98_fu_9574_p2 = (b_251_fu_9569_p2 & a_312_fu_9563_p2);

assign z1_99_fu_9655_p2 = (b_255_fu_9650_p2 & a_316_fu_9644_p2);

assign z1_9_fu_1278_p2 = (b_31_fu_1272_p2 & a_37_fu_1266_p2);

assign z1_fu_598_p2 = (b_5_fu_592_p2 & a_9_fu_586_p2);

assign z2_100_fu_9715_p2 = (b1_168_reg_14473_pp0_iter1_reg & a1_375_fu_9686_p3);

assign z2_102_fu_9820_p2 = (a1_377_fu_9796_p3 & a1_309_reg_14069_pp0_iter1_reg);

assign z2_103_fu_9900_p2 = (b1_170_reg_14479_pp0_iter1_reg & a1_378_fu_9865_p3);

assign z2_104_fu_9949_p2 = (a1_379_fu_9925_p3 & a1_310_reg_14085_pp0_iter1_reg);

assign z2_107_fu_10197_p2 = (b1_173_reg_14485_pp0_iter1_reg & a1_383_fu_10162_p3);

assign z2_108_fu_10278_p2 = (b1_174_reg_14498_pp0_iter1_reg & a1_384_fu_10242_p3);

assign z2_109_fu_10332_p2 = (b1_175_reg_14504_pp0_iter1_reg & a1_385_fu_10303_p3);

assign z2_10_fu_1456_p2 = (b1_109_fu_1424_p3 & a1_275_fu_1416_p3);

assign z2_111_fu_10485_p2 = (b1_177_reg_14518_pp0_iter1_reg & a1_387_fu_10449_p3);

assign z2_112_fu_10566_p2 = (b1_178_reg_14531_pp0_iter1_reg & a1_388_fu_10530_p3);

assign z2_113_fu_10620_p2 = (b1_179_reg_14537_pp0_iter1_reg & a1_389_fu_10591_p3);

assign z2_115_fu_10730_p2 = (b1_181_reg_14543_pp0_iter1_reg & a1_391_fu_10701_p3);

assign z2_116_fu_10810_p2 = (b1_182_reg_14556_pp0_iter1_reg & a1_392_fu_10775_p3);

assign z2_117_fu_10864_p2 = (b1_183_reg_14562_pp0_iter1_reg & a1_393_fu_10835_p3);

assign z2_120_fu_11041_p2 = (a1_397_fu_11017_p3 & a1_311_reg_14095_pp0_iter1_reg);

assign z2_121_fu_11121_p2 = (b1_185_reg_14568_pp0_iter1_reg & a1_398_fu_11086_p3);

assign z2_122_fu_11170_p2 = (a1_399_fu_11146_p3 & a1_312_reg_14111_pp0_iter1_reg);

assign z2_124_fu_11308_p2 = (b1_187_reg_14574_pp0_iter1_reg & a1_401_fu_11273_p3);

assign z2_125_fu_11389_p2 = (b1_188_reg_14587_pp0_iter1_reg & a1_402_fu_11353_p3);

assign z2_126_fu_11443_p2 = (b1_189_reg_14593_pp0_iter1_reg & a1_403_fu_11414_p3);

assign z2_128_fu_11548_p2 = (a1_405_fu_11524_p3 & a1_313_reg_14128_pp0_iter1_reg);

assign z2_129_fu_11628_p2 = (b1_190_reg_14599_pp0_iter1_reg & a1_406_fu_11593_p3);

assign z2_130_fu_11677_p2 = (a1_407_fu_11653_p3 & a1_261_reg_13605_pp0_iter1_reg);

assign z2_134_fu_11926_p2 = (b1_99_reg_13628_pp0_iter1_reg & a1_369_fu_9291_p3);

assign z2_135_fu_11961_p2 = (b1_100_reg_13648_pp0_iter1_reg & a1_370_fu_9360_p3);

assign z2_136_fu_11996_p2 = (b1_101_reg_13658_pp0_iter1_reg & a1_371_fu_9420_p3);

assign z2_138_fu_12077_p2 = (b1_103_reg_13678_pp0_iter1_reg & a1_373_fu_9545_p3);

assign z2_139_fu_12112_p2 = (b1_104_reg_13698_pp0_iter1_reg & a1_374_fu_9625_p3);

assign z2_13_fu_1840_p2 = (b1_112_fu_1808_p3 & a1_279_fu_1794_p3);

assign z2_140_fu_12147_p2 = (b1_105_reg_13708_pp0_iter1_reg & a1_375_fu_9686_p3);

assign z2_142_fu_12228_p2 = (b1_107_reg_13718_pp0_iter1_reg & a1_377_fu_9796_p3);

assign z2_143_fu_12263_p2 = (b1_108_reg_13738_pp0_iter1_reg & a1_378_fu_9865_p3);

assign z2_144_fu_12298_p2 = (b1_109_reg_13748_pp0_iter1_reg & a1_379_fu_9925_p3);

assign z2_147_fu_12451_p2 = (b1_112_reg_13768_pp0_iter1_reg & a1_383_fu_10162_p3);

assign z2_148_fu_12486_p2 = (b1_113_reg_13788_pp0_iter1_reg & a1_384_fu_10242_p3);

assign z2_149_fu_12521_p2 = (b1_114_reg_13798_pp0_iter1_reg & a1_385_fu_10303_p3);

assign z2_14_fu_1946_p2 = (b1_113_fu_1914_p3 & a1_280_fu_1900_p3);

assign z2_151_fu_12602_p2 = (b1_116_reg_13818_pp0_iter1_reg & a1_387_fu_10449_p3);

assign z2_152_fu_12637_p2 = (b1_117_reg_13838_pp0_iter1_reg & a1_388_fu_10530_p3);

assign z2_153_fu_12672_p2 = (b1_118_reg_13848_pp0_iter1_reg & a1_389_fu_10591_p3);

assign z2_155_fu_12753_p2 = (b1_120_reg_13858_pp0_iter1_reg & a1_391_fu_10701_p3);

assign z2_156_fu_12788_p2 = (b1_121_reg_13878_pp0_iter1_reg & a1_392_fu_10775_p3);

assign z2_157_fu_12823_p2 = (b1_122_reg_13888_pp0_iter1_reg & a1_393_fu_10835_p3);

assign z2_15_fu_2012_p2 = (b1_114_fu_1980_p3 & a1_281_fu_1972_p3);

assign z2_160_fu_12976_p2 = (b1_125_reg_13898_pp0_iter1_reg & a1_397_fu_11017_p3);

assign z2_161_fu_13011_p2 = (b1_126_reg_13918_pp0_iter1_reg & a1_398_fu_11086_p3);

assign z2_162_fu_13046_p2 = (b1_127_reg_13928_pp0_iter1_reg & a1_399_fu_11146_p3);

assign z2_164_fu_13127_p2 = (b1_129_reg_13948_pp0_iter1_reg & a1_401_fu_11273_p3);

assign z2_165_fu_13162_p2 = (b1_130_reg_13968_pp0_iter1_reg & a1_402_fu_11353_p3);

assign z2_166_fu_13197_p2 = (b1_131_reg_13978_pp0_iter1_reg & a1_403_fu_11414_p3);

assign z2_168_fu_13278_p2 = (b1_133_reg_13988_pp0_iter1_reg & a1_405_fu_11524_p3);

assign z2_169_fu_13313_p2 = (b1_134_reg_14008_pp0_iter1_reg & a1_406_fu_11593_p3);

assign z2_170_fu_13348_p2 = (b1_135_reg_14018_pp0_iter1_reg & a1_407_fu_11653_p3);

assign z2_174_fu_794_p3 = {{a1_13_fu_782_p2}, {a0_fu_788_p2}};

assign z2_175_fu_1170_p3 = {{a1_19_fu_1158_p2}, {a0_16_fu_1164_p2}};

assign z2_176_fu_1474_p3 = {{a1_24_fu_1462_p2}, {a0_23_fu_1468_p2}};

assign z2_177_fu_1520_p3 = {{a1_276_fu_1508_p2}, {a0_24_fu_1514_p2}};

assign z2_178_fu_2030_p3 = {{a1_34_fu_2018_p2}, {a0_36_fu_2024_p2}};

assign z2_179_fu_2406_p3 = {{a1_40_fu_2394_p2}, {a0_45_fu_2400_p2}};

assign z2_17_fu_2216_p2 = (b1_116_fu_2184_p3 & a1_283_fu_2170_p3);

assign z2_180_fu_2710_p3 = {{a1_46_fu_2698_p2}, {a0_49_fu_2704_p2}};

assign z2_181_fu_2756_p3 = {{a1_290_fu_2744_p2}, {a0_50_fu_2750_p2}};

assign z2_182_fu_3130_p3 = {{a1_56_fu_3118_p2}, {a0_57_fu_3124_p2}};

assign z2_183_fu_3506_p3 = {{a1_61_fu_3494_p2}, {a0_64_fu_3500_p2}};

assign z2_184_fu_3810_p3 = {{a1_66_fu_3798_p2}, {a0_69_fu_3804_p2}};

assign z2_185_fu_3856_p3 = {{a1_304_fu_3844_p2}, {a0_70_fu_3850_p2}};

assign z2_186_fu_3952_p3 = {{a1_305_fu_3928_p2}, {a0_73_fu_3934_p2}};

assign z2_187_fu_6098_p3 = {{a1_98_fu_6086_p2}, {a0_111_fu_6092_p2}};

assign z2_188_fu_6296_p3 = {{a1_103_fu_6284_p2}, {a0_117_fu_6290_p2}};

assign z2_189_fu_6480_p3 = {{a1_109_fu_6468_p2}, {a0_128_fu_6474_p2}};

assign z2_18_fu_2322_p2 = (b1_117_fu_2290_p3 & a1_284_fu_2276_p3);

assign z2_190_fu_6526_p3 = {{a1_332_fu_6514_p2}, {a0_129_fu_6520_p2}};

assign z2_191_fu_7140_p3 = {{a1_126_fu_7128_p2}, {a0_150_fu_7134_p2}};

assign z2_192_fu_7716_p3 = {{a1_141_fu_7704_p2}, {a0_167_fu_7710_p2}};

assign z2_193_fu_7853_p3 = {{a1_142_fu_7841_p2}, {a0_170_fu_7847_p2}};

assign z2_194_fu_8075_p3 = {{a1_149_fu_8063_p2}, {a0_190_fu_8069_p2}};

assign z2_195_fu_8348_p3 = {{a1_155_fu_8336_p2}, {a0_195_fu_8342_p2}};

assign z2_196_fu_8568_p3 = {{a1_161_fu_8556_p2}, {a0_200_fu_8562_p2}};

assign z2_197_fu_8614_p3 = {{a1_364_fu_8602_p2}, {a0_201_fu_8608_p2}};

assign z2_198_fu_8795_p3 = {{a1_164_fu_8783_p2}, {a0_203_fu_8789_p2}};

assign z2_199_fu_8946_p3 = {{a1_165_fu_8934_p2}, {a0_204_fu_8940_p2}};

assign z2_19_fu_2388_p2 = (b1_118_fu_2356_p3 & a1_285_fu_2348_p3);

assign z2_1_fu_710_p2 = (b1_100_fu_678_p3 & a1_266_fu_664_p3);

assign z2_200_fu_9097_p3 = {{a1_167_fu_9085_p2}, {a0_205_fu_9091_p2}};

assign z2_201_fu_9143_p3 = {{a1_365_fu_9131_p2}, {a0_206_fu_9137_p2}};

assign z2_202_fu_9461_p3 = {{a1_178_fu_9449_p2}, {a0_214_fu_9455_p2}};

assign z2_203_fu_9732_p3 = {{a1_183_fu_9720_p2}, {a0_219_fu_9726_p2}};

assign z2_204_fu_9966_p3 = {{a1_190_fu_9954_p2}, {a0_224_fu_9960_p2}};

assign z2_205_fu_10012_p3 = {{a1_380_fu_10000_p2}, {a0_225_fu_10006_p2}};

assign z2_206_fu_10349_p3 = {{a1_198_fu_10337_p2}, {a0_232_fu_10343_p2}};

assign z2_207_fu_10637_p3 = {{a1_212_fu_10625_p2}, {a0_237_fu_10631_p2}};

assign z2_208_fu_10881_p3 = {{a1_217_fu_10869_p2}, {a0_242_fu_10875_p2}};

assign z2_209_fu_10927_p3 = {{a1_394_fu_10915_p2}, {a0_243_fu_10921_p2}};

assign z2_210_fu_11187_p3 = {{a1_225_fu_11175_p2}, {a0_250_fu_11181_p2}};

assign z2_211_fu_11460_p3 = {{a1_230_fu_11448_p2}, {a0_255_fu_11454_p2}};

assign z2_212_fu_11694_p3 = {{a1_fu_11682_p2}, {a0_260_fu_11688_p2}};

assign z2_213_fu_11740_p3 = {{a1_408_fu_11728_p2}, {a0_261_fu_11734_p2}};

assign z2_214_fu_11812_p3 = {{a1_409_fu_11800_p2}, {a0_263_fu_11806_p2}};

assign z2_215_fu_12013_p3 = {{a1_240_fu_12001_p2}, {a0_266_fu_12007_p2}};

assign z2_216_fu_12164_p3 = {{a1_241_fu_12152_p2}, {a0_267_fu_12158_p2}};

assign z2_217_fu_12315_p3 = {{a1_242_fu_12303_p2}, {a0_268_fu_12309_p2}};

assign z2_218_fu_12361_p3 = {{a1_411_fu_12349_p2}, {a0_269_fu_12355_p2}};

assign z2_219_fu_12538_p3 = {{a1_245_fu_12526_p2}, {a0_271_fu_12532_p2}};

assign z2_21_fu_2520_p2 = (b1_120_fu_2488_p3 & a1_287_fu_2480_p3);

assign z2_220_fu_12689_p3 = {{a1_246_fu_12677_p2}, {a0_272_fu_12683_p2}};

assign z2_221_fu_12840_p3 = {{a1_247_fu_12828_p2}, {a0_273_fu_12834_p2}};

assign z2_222_fu_12886_p3 = {{a1_412_fu_12874_p2}, {a0_274_fu_12880_p2}};

assign z2_223_fu_13063_p3 = {{a1_250_fu_13051_p2}, {a0_276_fu_13057_p2}};

assign z2_224_fu_13214_p3 = {{a1_251_fu_13202_p2}, {a0_277_fu_13208_p2}};

assign z2_225_fu_13365_p3 = {{a1_252_fu_13353_p2}, {a0_278_fu_13359_p2}};

assign z2_226_fu_13411_p3 = {{a1_413_fu_13399_p2}, {a0_279_fu_13405_p2}};

assign z2_227_fu_13483_p3 = {{a1_414_fu_13471_p2}, {a0_281_fu_13477_p2}};

assign z2_22_fu_2626_p2 = (b1_121_fu_2594_p3 & a1_288_fu_2580_p3);

assign z2_23_fu_2692_p2 = (b1_122_fu_2660_p3 & a1_289_fu_2652_p3);

assign z2_26_fu_2940_p2 = (b1_125_fu_2908_p3 & a1_293_fu_2900_p3);

assign z2_27_fu_3046_p2 = (b1_126_fu_3014_p3 & a1_294_fu_3000_p3);

assign z2_28_fu_3112_p2 = (b1_127_fu_3080_p3 & a1_295_fu_3072_p3);

assign z2_2_fu_776_p2 = (b1_101_fu_744_p3 & a1_267_fu_736_p3);

assign z2_30_fu_3316_p2 = (b1_129_fu_3284_p3 & a1_297_fu_3270_p3);

assign z2_31_fu_3422_p2 = (b1_130_fu_3390_p3 & a1_298_fu_3376_p3);

assign z2_32_fu_3488_p2 = (b1_131_fu_3456_p3 & a1_299_fu_3448_p3);

assign z2_34_fu_3620_p2 = (b1_133_fu_3588_p3 & a1_301_fu_3580_p3);

assign z2_35_fu_3726_p2 = (b1_134_fu_3694_p3 & a1_302_fu_3680_p3);

assign z2_36_fu_3792_p2 = (b1_135_fu_3760_p3 & a1_303_fu_3752_p3);

assign z2_40_fu_5986_p2 = (b1_138_reg_14190 & a1_321_reg_14175);

assign z2_41_fu_6040_p2 = (b1_139_reg_14218 & a1_322_reg_14212);

assign z2_42_fu_6082_p2 = (b1_140_reg_14231 & a1_323_reg_14225);

assign z2_44_fu_6182_p2 = (b1_142_reg_14261 & a1_325_reg_14255);

assign z2_45_fu_6238_p2 = (b1_143_reg_14289 & a1_326_reg_14283);

assign z2_46_fu_6280_p2 = (b1_144_reg_14302 & a1_327_reg_14296);

assign z2_48_fu_6368_p2 = (b1_146_reg_14315 & a1_329_reg_14309);

assign z2_49_fu_6422_p2 = (b1_147_reg_14343 & a1_330_reg_14337);

assign z2_4_fu_980_p2 = (b1_103_fu_948_p3 & a1_269_fu_934_p3);

assign z2_50_fu_6464_p2 = (b1_148_reg_14356 & a1_331_reg_14350);

assign z2_53_fu_6950_p2 = (b1_150_fu_6918_p3 & a1_339_fu_6904_p3);

assign z2_54_fu_7056_p2 = (b1_151_fu_7024_p3 & a1_340_fu_7010_p3);

assign z2_55_fu_7122_p2 = (b1_152_fu_7090_p3 & a1_341_fu_7082_p3);

assign z2_57_fu_7402_p2 = (b1_153_fu_7370_p3 & a1_344_fu_7362_p3);

assign z2_58_fu_7504_p2 = (a1_346_fu_7474_p2 & a1_343_fu_7328_p3);

assign z2_59_fu_7534_p2 = (b1_153_fu_7370_p3 & a1_346_fu_7474_p2);

assign z2_5_fu_1086_p2 = (b1_104_fu_1054_p3 & a1_270_fu_1040_p3);

assign z2_60_fu_7598_p2 = (a1_348_reg_14777 & a1_342_reg_14752);

assign z2_61_fu_7667_p2 = (b1_154_reg_14798 & a1_349_fu_7632_p3);

assign z2_62_fu_7700_p2 = (a1_350_reg_14762 & a1_337_reg_14691);

assign z2_64_fu_7770_p2 = (b1_150_reg_14706 & a1_348_reg_14777);

assign z2_65_fu_7804_p2 = (b1_151_reg_14726 & a1_349_fu_7632_p3);

assign z2_66_fu_7837_p2 = (b1_152_reg_14736 & a1_350_reg_14762);

assign z2_68_fu_7939_p2 = (a1_353_fu_7915_p3 & a1_333_reg_14371_pp0_iter1_reg);

assign z2_69_fu_8009_p2 = (b1_156_reg_14411_pp0_iter1_reg & a1_354_fu_7974_p3);

assign z2_6_fu_1152_p2 = (b1_105_fu_1120_p3 & a1_271_fu_1112_p3);

assign z2_70_fu_8058_p2 = (a1_355_fu_8034_p3 & a1_334_reg_14385_pp0_iter1_reg);

assign z2_72_fu_8196_p2 = (b1_158_reg_14417_pp0_iter1_reg & a1_357_fu_8161_p3);

assign z2_73_fu_8277_p2 = (b1_159_reg_14430_pp0_iter1_reg & a1_358_fu_8241_p3);

assign z2_74_fu_8331_p2 = (b1_160_reg_14436_pp0_iter1_reg & a1_359_fu_8302_p3);

assign z2_76_fu_8426_p2 = (a1_361_fu_8402_p3 & a1_335_reg_14397_pp0_iter1_reg);

assign z2_77_fu_8502_p2 = (b1_161_reg_14442_pp0_iter1_reg & a1_362_fu_8467_p3);

assign z2_78_fu_8551_p2 = (a1_363_fu_8527_p3 & a1_318_reg_14145_pp0_iter1_reg);

assign z2_81_fu_8708_p2 = (b1_138_reg_14190_pp0_iter1_reg & a1_353_fu_7915_p3);

assign z2_82_fu_8743_p2 = (b1_139_reg_14218_pp0_iter1_reg & a1_354_fu_7974_p3);

assign z2_83_fu_8778_p2 = (b1_140_reg_14231_pp0_iter1_reg & a1_355_fu_8034_p3);

assign z2_85_fu_8859_p2 = (b1_142_reg_14261_pp0_iter1_reg & a1_357_fu_8161_p3);

assign z2_86_fu_8894_p2 = (b1_143_reg_14289_pp0_iter1_reg & a1_358_fu_8241_p3);

assign z2_87_fu_8929_p2 = (b1_144_reg_14302_pp0_iter1_reg & a1_359_fu_8302_p3);

assign z2_89_fu_9010_p2 = (b1_146_reg_14315_pp0_iter1_reg & a1_361_fu_8402_p3);

assign z2_8_fu_1284_p2 = (b1_107_fu_1252_p3 & a1_273_fu_1244_p3);

assign z2_90_fu_9045_p2 = (b1_147_reg_14343_pp0_iter1_reg & a1_362_fu_8467_p3);

assign z2_91_fu_9080_p2 = (b1_148_reg_14356_pp0_iter1_reg & a1_363_fu_8527_p3);

assign z2_94_fu_9315_p2 = (a1_369_fu_9291_p3 & a1_307_reg_14036_pp0_iter1_reg);

assign z2_95_fu_9395_p2 = (b1_164_reg_14448_pp0_iter1_reg & a1_370_fu_9360_p3);

assign z2_96_fu_9444_p2 = (a1_371_fu_9420_p3 & a1_308_reg_14052_pp0_iter1_reg);

assign z2_98_fu_9580_p2 = (b1_166_reg_14454_pp0_iter1_reg & a1_373_fu_9545_p3);

assign z2_99_fu_9661_p2 = (b1_167_reg_14467_pp0_iter1_reg & a1_374_fu_9625_p3);

assign z2_9_fu_1390_p2 = (b1_108_fu_1358_p3 & a1_274_fu_1344_p3);

assign z2_fu_604_p2 = (b1_99_fu_572_p3 & a1_265_fu_558_p3);

endmodule //binary_tower_32b_inv
